module TensorLoadNarrowVME_1(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [7:0]   io_vme_rd_cmd_bits_len,
  output [20:0]  io_vme_rd_cmd_bits_tag,
  output         io_vme_rd_data_ready,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input  [20:0]  io_vme_rd_data_bits_tag,
  input          io_tensor_rd_0_idx_valid,
  input  [9:0]   io_tensor_rd_0_idx_bits,
  output         io_tensor_rd_0_data_valid,
  output [31:0]  io_tensor_rd_0_data_bits_0_0,
  output [31:0]  io_tensor_rd_0_data_bits_0_1,
  output [31:0]  io_tensor_rd_0_data_bits_0_2,
  output [31:0]  io_tensor_rd_0_data_bits_0_3,
  output [31:0]  io_tensor_rd_0_data_bits_0_4,
  output [31:0]  io_tensor_rd_0_data_bits_0_5,
  output [31:0]  io_tensor_rd_0_data_bits_0_6,
  output [31:0]  io_tensor_rd_0_data_bits_0_7,
  output [31:0]  io_tensor_rd_0_data_bits_0_8,
  output [31:0]  io_tensor_rd_0_data_bits_0_9,
  output [31:0]  io_tensor_rd_0_data_bits_0_10,
  output [31:0]  io_tensor_rd_0_data_bits_0_11,
  output [31:0]  io_tensor_rd_0_data_bits_0_12,
  output [31:0]  io_tensor_rd_0_data_bits_0_13,
  output [31:0]  io_tensor_rd_0_data_bits_0_14,
  output [31:0]  io_tensor_rd_0_data_bits_0_15,
  output [31:0]  io_tensor_rd_0_data_bits_1_0,
  output [31:0]  io_tensor_rd_0_data_bits_1_1,
  output [31:0]  io_tensor_rd_0_data_bits_1_2,
  output [31:0]  io_tensor_rd_0_data_bits_1_3,
  output [31:0]  io_tensor_rd_0_data_bits_1_4,
  output [31:0]  io_tensor_rd_0_data_bits_1_5,
  output [31:0]  io_tensor_rd_0_data_bits_1_6,
  output [31:0]  io_tensor_rd_0_data_bits_1_7,
  output [31:0]  io_tensor_rd_0_data_bits_1_8,
  output [31:0]  io_tensor_rd_0_data_bits_1_9,
  output [31:0]  io_tensor_rd_0_data_bits_1_10,
  output [31:0]  io_tensor_rd_0_data_bits_1_11,
  output [31:0]  io_tensor_rd_0_data_bits_1_12,
  output [31:0]  io_tensor_rd_0_data_bits_1_13,
  output [31:0]  io_tensor_rd_0_data_bits_1_14,
  output [31:0]  io_tensor_rd_0_data_bits_1_15,
  output [31:0]  io_tensor_rd_0_data_bits_2_0,
  output [31:0]  io_tensor_rd_0_data_bits_2_1,
  output [31:0]  io_tensor_rd_0_data_bits_2_2,
  output [31:0]  io_tensor_rd_0_data_bits_2_3,
  output [31:0]  io_tensor_rd_0_data_bits_2_4,
  output [31:0]  io_tensor_rd_0_data_bits_2_5,
  output [31:0]  io_tensor_rd_0_data_bits_2_6,
  output [31:0]  io_tensor_rd_0_data_bits_2_7,
  output [31:0]  io_tensor_rd_0_data_bits_2_8,
  output [31:0]  io_tensor_rd_0_data_bits_2_9,
  output [31:0]  io_tensor_rd_0_data_bits_2_10,
  output [31:0]  io_tensor_rd_0_data_bits_2_11,
  output [31:0]  io_tensor_rd_0_data_bits_2_12,
  output [31:0]  io_tensor_rd_0_data_bits_2_13,
  output [31:0]  io_tensor_rd_0_data_bits_2_14,
  output [31:0]  io_tensor_rd_0_data_bits_2_15,
  output [31:0]  io_tensor_rd_0_data_bits_3_0,
  output [31:0]  io_tensor_rd_0_data_bits_3_1,
  output [31:0]  io_tensor_rd_0_data_bits_3_2,
  output [31:0]  io_tensor_rd_0_data_bits_3_3,
  output [31:0]  io_tensor_rd_0_data_bits_3_4,
  output [31:0]  io_tensor_rd_0_data_bits_3_5,
  output [31:0]  io_tensor_rd_0_data_bits_3_6,
  output [31:0]  io_tensor_rd_0_data_bits_3_7,
  output [31:0]  io_tensor_rd_0_data_bits_3_8,
  output [31:0]  io_tensor_rd_0_data_bits_3_9,
  output [31:0]  io_tensor_rd_0_data_bits_3_10,
  output [31:0]  io_tensor_rd_0_data_bits_3_11,
  output [31:0]  io_tensor_rd_0_data_bits_3_12,
  output [31:0]  io_tensor_rd_0_data_bits_3_13,
  output [31:0]  io_tensor_rd_0_data_bits_3_14,
  output [31:0]  io_tensor_rd_0_data_bits_3_15,
  output [31:0]  io_tensor_rd_0_data_bits_4_0,
  output [31:0]  io_tensor_rd_0_data_bits_4_1,
  output [31:0]  io_tensor_rd_0_data_bits_4_2,
  output [31:0]  io_tensor_rd_0_data_bits_4_3,
  output [31:0]  io_tensor_rd_0_data_bits_4_4,
  output [31:0]  io_tensor_rd_0_data_bits_4_5,
  output [31:0]  io_tensor_rd_0_data_bits_4_6,
  output [31:0]  io_tensor_rd_0_data_bits_4_7,
  output [31:0]  io_tensor_rd_0_data_bits_4_8,
  output [31:0]  io_tensor_rd_0_data_bits_4_9,
  output [31:0]  io_tensor_rd_0_data_bits_4_10,
  output [31:0]  io_tensor_rd_0_data_bits_4_11,
  output [31:0]  io_tensor_rd_0_data_bits_4_12,
  output [31:0]  io_tensor_rd_0_data_bits_4_13,
  output [31:0]  io_tensor_rd_0_data_bits_4_14,
  output [31:0]  io_tensor_rd_0_data_bits_4_15,
  output [31:0]  io_tensor_rd_0_data_bits_5_0,
  output [31:0]  io_tensor_rd_0_data_bits_5_1,
  output [31:0]  io_tensor_rd_0_data_bits_5_2,
  output [31:0]  io_tensor_rd_0_data_bits_5_3,
  output [31:0]  io_tensor_rd_0_data_bits_5_4,
  output [31:0]  io_tensor_rd_0_data_bits_5_5,
  output [31:0]  io_tensor_rd_0_data_bits_5_6,
  output [31:0]  io_tensor_rd_0_data_bits_5_7,
  output [31:0]  io_tensor_rd_0_data_bits_5_8,
  output [31:0]  io_tensor_rd_0_data_bits_5_9,
  output [31:0]  io_tensor_rd_0_data_bits_5_10,
  output [31:0]  io_tensor_rd_0_data_bits_5_11,
  output [31:0]  io_tensor_rd_0_data_bits_5_12,
  output [31:0]  io_tensor_rd_0_data_bits_5_13,
  output [31:0]  io_tensor_rd_0_data_bits_5_14,
  output [31:0]  io_tensor_rd_0_data_bits_5_15,
  output [31:0]  io_tensor_rd_0_data_bits_6_0,
  output [31:0]  io_tensor_rd_0_data_bits_6_1,
  output [31:0]  io_tensor_rd_0_data_bits_6_2,
  output [31:0]  io_tensor_rd_0_data_bits_6_3,
  output [31:0]  io_tensor_rd_0_data_bits_6_4,
  output [31:0]  io_tensor_rd_0_data_bits_6_5,
  output [31:0]  io_tensor_rd_0_data_bits_6_6,
  output [31:0]  io_tensor_rd_0_data_bits_6_7,
  output [31:0]  io_tensor_rd_0_data_bits_6_8,
  output [31:0]  io_tensor_rd_0_data_bits_6_9,
  output [31:0]  io_tensor_rd_0_data_bits_6_10,
  output [31:0]  io_tensor_rd_0_data_bits_6_11,
  output [31:0]  io_tensor_rd_0_data_bits_6_12,
  output [31:0]  io_tensor_rd_0_data_bits_6_13,
  output [31:0]  io_tensor_rd_0_data_bits_6_14,
  output [31:0]  io_tensor_rd_0_data_bits_6_15,
  output [31:0]  io_tensor_rd_0_data_bits_7_0,
  output [31:0]  io_tensor_rd_0_data_bits_7_1,
  output [31:0]  io_tensor_rd_0_data_bits_7_2,
  output [31:0]  io_tensor_rd_0_data_bits_7_3,
  output [31:0]  io_tensor_rd_0_data_bits_7_4,
  output [31:0]  io_tensor_rd_0_data_bits_7_5,
  output [31:0]  io_tensor_rd_0_data_bits_7_6,
  output [31:0]  io_tensor_rd_0_data_bits_7_7,
  output [31:0]  io_tensor_rd_0_data_bits_7_8,
  output [31:0]  io_tensor_rd_0_data_bits_7_9,
  output [31:0]  io_tensor_rd_0_data_bits_7_10,
  output [31:0]  io_tensor_rd_0_data_bits_7_11,
  output [31:0]  io_tensor_rd_0_data_bits_7_12,
  output [31:0]  io_tensor_rd_0_data_bits_7_13,
  output [31:0]  io_tensor_rd_0_data_bits_7_14,
  output [31:0]  io_tensor_rd_0_data_bits_7_15,
  output [31:0]  io_tensor_rd_0_data_bits_8_0,
  output [31:0]  io_tensor_rd_0_data_bits_8_1,
  output [31:0]  io_tensor_rd_0_data_bits_8_2,
  output [31:0]  io_tensor_rd_0_data_bits_8_3,
  output [31:0]  io_tensor_rd_0_data_bits_8_4,
  output [31:0]  io_tensor_rd_0_data_bits_8_5,
  output [31:0]  io_tensor_rd_0_data_bits_8_6,
  output [31:0]  io_tensor_rd_0_data_bits_8_7,
  output [31:0]  io_tensor_rd_0_data_bits_8_8,
  output [31:0]  io_tensor_rd_0_data_bits_8_9,
  output [31:0]  io_tensor_rd_0_data_bits_8_10,
  output [31:0]  io_tensor_rd_0_data_bits_8_11,
  output [31:0]  io_tensor_rd_0_data_bits_8_12,
  output [31:0]  io_tensor_rd_0_data_bits_8_13,
  output [31:0]  io_tensor_rd_0_data_bits_8_14,
  output [31:0]  io_tensor_rd_0_data_bits_8_15,
  output [31:0]  io_tensor_rd_0_data_bits_9_0,
  output [31:0]  io_tensor_rd_0_data_bits_9_1,
  output [31:0]  io_tensor_rd_0_data_bits_9_2,
  output [31:0]  io_tensor_rd_0_data_bits_9_3,
  output [31:0]  io_tensor_rd_0_data_bits_9_4,
  output [31:0]  io_tensor_rd_0_data_bits_9_5,
  output [31:0]  io_tensor_rd_0_data_bits_9_6,
  output [31:0]  io_tensor_rd_0_data_bits_9_7,
  output [31:0]  io_tensor_rd_0_data_bits_9_8,
  output [31:0]  io_tensor_rd_0_data_bits_9_9,
  output [31:0]  io_tensor_rd_0_data_bits_9_10,
  output [31:0]  io_tensor_rd_0_data_bits_9_11,
  output [31:0]  io_tensor_rd_0_data_bits_9_12,
  output [31:0]  io_tensor_rd_0_data_bits_9_13,
  output [31:0]  io_tensor_rd_0_data_bits_9_14,
  output [31:0]  io_tensor_rd_0_data_bits_9_15,
  output [31:0]  io_tensor_rd_0_data_bits_10_0,
  output [31:0]  io_tensor_rd_0_data_bits_10_1,
  output [31:0]  io_tensor_rd_0_data_bits_10_2,
  output [31:0]  io_tensor_rd_0_data_bits_10_3,
  output [31:0]  io_tensor_rd_0_data_bits_10_4,
  output [31:0]  io_tensor_rd_0_data_bits_10_5,
  output [31:0]  io_tensor_rd_0_data_bits_10_6,
  output [31:0]  io_tensor_rd_0_data_bits_10_7,
  output [31:0]  io_tensor_rd_0_data_bits_10_8,
  output [31:0]  io_tensor_rd_0_data_bits_10_9,
  output [31:0]  io_tensor_rd_0_data_bits_10_10,
  output [31:0]  io_tensor_rd_0_data_bits_10_11,
  output [31:0]  io_tensor_rd_0_data_bits_10_12,
  output [31:0]  io_tensor_rd_0_data_bits_10_13,
  output [31:0]  io_tensor_rd_0_data_bits_10_14,
  output [31:0]  io_tensor_rd_0_data_bits_10_15,
  output [31:0]  io_tensor_rd_0_data_bits_11_0,
  output [31:0]  io_tensor_rd_0_data_bits_11_1,
  output [31:0]  io_tensor_rd_0_data_bits_11_2,
  output [31:0]  io_tensor_rd_0_data_bits_11_3,
  output [31:0]  io_tensor_rd_0_data_bits_11_4,
  output [31:0]  io_tensor_rd_0_data_bits_11_5,
  output [31:0]  io_tensor_rd_0_data_bits_11_6,
  output [31:0]  io_tensor_rd_0_data_bits_11_7,
  output [31:0]  io_tensor_rd_0_data_bits_11_8,
  output [31:0]  io_tensor_rd_0_data_bits_11_9,
  output [31:0]  io_tensor_rd_0_data_bits_11_10,
  output [31:0]  io_tensor_rd_0_data_bits_11_11,
  output [31:0]  io_tensor_rd_0_data_bits_11_12,
  output [31:0]  io_tensor_rd_0_data_bits_11_13,
  output [31:0]  io_tensor_rd_0_data_bits_11_14,
  output [31:0]  io_tensor_rd_0_data_bits_11_15,
  output [31:0]  io_tensor_rd_0_data_bits_12_0,
  output [31:0]  io_tensor_rd_0_data_bits_12_1,
  output [31:0]  io_tensor_rd_0_data_bits_12_2,
  output [31:0]  io_tensor_rd_0_data_bits_12_3,
  output [31:0]  io_tensor_rd_0_data_bits_12_4,
  output [31:0]  io_tensor_rd_0_data_bits_12_5,
  output [31:0]  io_tensor_rd_0_data_bits_12_6,
  output [31:0]  io_tensor_rd_0_data_bits_12_7,
  output [31:0]  io_tensor_rd_0_data_bits_12_8,
  output [31:0]  io_tensor_rd_0_data_bits_12_9,
  output [31:0]  io_tensor_rd_0_data_bits_12_10,
  output [31:0]  io_tensor_rd_0_data_bits_12_11,
  output [31:0]  io_tensor_rd_0_data_bits_12_12,
  output [31:0]  io_tensor_rd_0_data_bits_12_13,
  output [31:0]  io_tensor_rd_0_data_bits_12_14,
  output [31:0]  io_tensor_rd_0_data_bits_12_15,
  output [31:0]  io_tensor_rd_0_data_bits_13_0,
  output [31:0]  io_tensor_rd_0_data_bits_13_1,
  output [31:0]  io_tensor_rd_0_data_bits_13_2,
  output [31:0]  io_tensor_rd_0_data_bits_13_3,
  output [31:0]  io_tensor_rd_0_data_bits_13_4,
  output [31:0]  io_tensor_rd_0_data_bits_13_5,
  output [31:0]  io_tensor_rd_0_data_bits_13_6,
  output [31:0]  io_tensor_rd_0_data_bits_13_7,
  output [31:0]  io_tensor_rd_0_data_bits_13_8,
  output [31:0]  io_tensor_rd_0_data_bits_13_9,
  output [31:0]  io_tensor_rd_0_data_bits_13_10,
  output [31:0]  io_tensor_rd_0_data_bits_13_11,
  output [31:0]  io_tensor_rd_0_data_bits_13_12,
  output [31:0]  io_tensor_rd_0_data_bits_13_13,
  output [31:0]  io_tensor_rd_0_data_bits_13_14,
  output [31:0]  io_tensor_rd_0_data_bits_13_15,
  output [31:0]  io_tensor_rd_0_data_bits_14_0,
  output [31:0]  io_tensor_rd_0_data_bits_14_1,
  output [31:0]  io_tensor_rd_0_data_bits_14_2,
  output [31:0]  io_tensor_rd_0_data_bits_14_3,
  output [31:0]  io_tensor_rd_0_data_bits_14_4,
  output [31:0]  io_tensor_rd_0_data_bits_14_5,
  output [31:0]  io_tensor_rd_0_data_bits_14_6,
  output [31:0]  io_tensor_rd_0_data_bits_14_7,
  output [31:0]  io_tensor_rd_0_data_bits_14_8,
  output [31:0]  io_tensor_rd_0_data_bits_14_9,
  output [31:0]  io_tensor_rd_0_data_bits_14_10,
  output [31:0]  io_tensor_rd_0_data_bits_14_11,
  output [31:0]  io_tensor_rd_0_data_bits_14_12,
  output [31:0]  io_tensor_rd_0_data_bits_14_13,
  output [31:0]  io_tensor_rd_0_data_bits_14_14,
  output [31:0]  io_tensor_rd_0_data_bits_14_15,
  output [31:0]  io_tensor_rd_0_data_bits_15_0,
  output [31:0]  io_tensor_rd_0_data_bits_15_1,
  output [31:0]  io_tensor_rd_0_data_bits_15_2,
  output [31:0]  io_tensor_rd_0_data_bits_15_3,
  output [31:0]  io_tensor_rd_0_data_bits_15_4,
  output [31:0]  io_tensor_rd_0_data_bits_15_5,
  output [31:0]  io_tensor_rd_0_data_bits_15_6,
  output [31:0]  io_tensor_rd_0_data_bits_15_7,
  output [31:0]  io_tensor_rd_0_data_bits_15_8,
  output [31:0]  io_tensor_rd_0_data_bits_15_9,
  output [31:0]  io_tensor_rd_0_data_bits_15_10,
  output [31:0]  io_tensor_rd_0_data_bits_15_11,
  output [31:0]  io_tensor_rd_0_data_bits_15_12,
  output [31:0]  io_tensor_rd_0_data_bits_15_13,
  output [31:0]  io_tensor_rd_0_data_bits_15_14,
  output [31:0]  io_tensor_rd_0_data_bits_15_15
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_255;
  reg [63:0] _RAND_258;
  reg [63:0] _RAND_261;
  reg [63:0] _RAND_264;
  reg [63:0] _RAND_267;
  reg [63:0] _RAND_270;
  reg [63:0] _RAND_273;
  reg [63:0] _RAND_276;
  reg [63:0] _RAND_279;
  reg [63:0] _RAND_282;
  reg [63:0] _RAND_285;
  reg [63:0] _RAND_288;
  reg [63:0] _RAND_291;
  reg [63:0] _RAND_294;
  reg [63:0] _RAND_297;
  reg [63:0] _RAND_300;
  reg [63:0] _RAND_303;
  reg [63:0] _RAND_306;
  reg [63:0] _RAND_309;
  reg [63:0] _RAND_312;
  reg [63:0] _RAND_315;
  reg [63:0] _RAND_318;
  reg [63:0] _RAND_321;
  reg [63:0] _RAND_324;
  reg [63:0] _RAND_327;
  reg [63:0] _RAND_330;
  reg [63:0] _RAND_333;
  reg [63:0] _RAND_336;
  reg [63:0] _RAND_339;
  reg [63:0] _RAND_342;
  reg [63:0] _RAND_345;
  reg [63:0] _RAND_348;
  reg [63:0] _RAND_351;
  reg [63:0] _RAND_354;
  reg [63:0] _RAND_357;
  reg [63:0] _RAND_360;
  reg [63:0] _RAND_363;
  reg [63:0] _RAND_366;
  reg [63:0] _RAND_369;
  reg [63:0] _RAND_372;
  reg [63:0] _RAND_375;
  reg [63:0] _RAND_378;
  reg [63:0] _RAND_381;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [63:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [127:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
`endif // RANDOMIZE_REG_INIT
  wire  vmeCmd_clock; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_reset; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_start; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_isBusy; // @[TensorLoadNarrowVME.scala 75:23]
  wire [127:0] vmeCmd_io_inst; // @[TensorLoadNarrowVME.scala 75:23]
  wire [31:0] vmeCmd_io_baddr; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_vmeCmd_ready; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_vmeCmd_valid; // @[TensorLoadNarrowVME.scala 75:23]
  wire [31:0] vmeCmd_io_vmeCmd_bits_addr; // @[TensorLoadNarrowVME.scala 75:23]
  wire [7:0] vmeCmd_io_vmeCmd_bits_len; // @[TensorLoadNarrowVME.scala 75:23]
  wire [20:0] vmeCmd_io_vmeCmd_bits_tag; // @[TensorLoadNarrowVME.scala 75:23]
  wire [8:0] vmeCmd_io_readLen; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_done; // @[TensorLoadNarrowVME.scala 75:23]
  wire  readData_clock; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_reset; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_start; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_vmeData_ready; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_vmeData_valid; // @[TensorLoadNarrowVME.scala 105:24]
  wire [20:0] readData_io_vmeData_bits_tag; // @[TensorLoadNarrowVME.scala 105:24]
  wire [9:0] readData_io_idx; // @[TensorLoadNarrowVME.scala 105:24]
  wire [6:0] readData_io_col; // @[TensorLoadNarrowVME.scala 105:24]
  wire  fillPadding_clock; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_reset; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_canWriteMem; // @[TensorLoadNarrowVME.scala 119:27]
  wire [127:0] fillPadding_io_inst; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_tensorIdx_valid; // @[TensorLoadNarrowVME.scala 119:27]
  wire [9:0] fillPadding_io_tensorIdx_bits; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_start; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_done; // @[TensorLoadNarrowVME.scala 119:27]
  reg [63:0] tensorFile_0 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_0_MPORT_128_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_0_MPORT_128_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_0_MPORT_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_0_MPORT_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_0_MPORT_128_en_pipe_0;
  reg [9:0] tensorFile_0_MPORT_128_addr_pipe_0;
  reg [63:0] tensorFile_1 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_1_MPORT_129_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_1_MPORT_129_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_1_MPORT_1_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_1_MPORT_1_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_1_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_1_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_1_MPORT_129_en_pipe_0;
  reg [9:0] tensorFile_1_MPORT_129_addr_pipe_0;
  reg [63:0] tensorFile_2 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_2_MPORT_130_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_2_MPORT_130_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_2_MPORT_2_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_2_MPORT_2_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_2_MPORT_2_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_2_MPORT_2_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_2_MPORT_130_en_pipe_0;
  reg [9:0] tensorFile_2_MPORT_130_addr_pipe_0;
  reg [63:0] tensorFile_3 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_3_MPORT_131_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_3_MPORT_131_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_3_MPORT_3_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_3_MPORT_3_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_3_MPORT_3_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_3_MPORT_3_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_3_MPORT_131_en_pipe_0;
  reg [9:0] tensorFile_3_MPORT_131_addr_pipe_0;
  reg [63:0] tensorFile_4 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_4_MPORT_132_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_4_MPORT_132_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_4_MPORT_4_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_4_MPORT_4_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_4_MPORT_4_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_4_MPORT_4_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_4_MPORT_132_en_pipe_0;
  reg [9:0] tensorFile_4_MPORT_132_addr_pipe_0;
  reg [63:0] tensorFile_5 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_5_MPORT_133_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_5_MPORT_133_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_5_MPORT_5_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_5_MPORT_5_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_5_MPORT_5_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_5_MPORT_5_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_5_MPORT_133_en_pipe_0;
  reg [9:0] tensorFile_5_MPORT_133_addr_pipe_0;
  reg [63:0] tensorFile_6 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_6_MPORT_134_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_6_MPORT_134_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_6_MPORT_6_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_6_MPORT_6_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_6_MPORT_6_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_6_MPORT_6_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_6_MPORT_134_en_pipe_0;
  reg [9:0] tensorFile_6_MPORT_134_addr_pipe_0;
  reg [63:0] tensorFile_7 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_7_MPORT_135_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_7_MPORT_135_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_7_MPORT_7_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_7_MPORT_7_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_7_MPORT_7_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_7_MPORT_7_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_7_MPORT_135_en_pipe_0;
  reg [9:0] tensorFile_7_MPORT_135_addr_pipe_0;
  reg [63:0] tensorFile_8 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_8_MPORT_136_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_8_MPORT_136_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_8_MPORT_8_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_8_MPORT_8_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_8_MPORT_8_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_8_MPORT_8_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_8_MPORT_136_en_pipe_0;
  reg [9:0] tensorFile_8_MPORT_136_addr_pipe_0;
  reg [63:0] tensorFile_9 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_9_MPORT_137_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_9_MPORT_137_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_9_MPORT_9_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_9_MPORT_9_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_9_MPORT_9_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_9_MPORT_9_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_9_MPORT_137_en_pipe_0;
  reg [9:0] tensorFile_9_MPORT_137_addr_pipe_0;
  reg [63:0] tensorFile_10 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_10_MPORT_138_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_10_MPORT_138_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_10_MPORT_10_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_10_MPORT_10_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_10_MPORT_10_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_10_MPORT_10_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_10_MPORT_138_en_pipe_0;
  reg [9:0] tensorFile_10_MPORT_138_addr_pipe_0;
  reg [63:0] tensorFile_11 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_11_MPORT_139_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_11_MPORT_139_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_11_MPORT_11_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_11_MPORT_11_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_11_MPORT_11_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_11_MPORT_11_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_11_MPORT_139_en_pipe_0;
  reg [9:0] tensorFile_11_MPORT_139_addr_pipe_0;
  reg [63:0] tensorFile_12 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_12_MPORT_140_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_12_MPORT_140_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_12_MPORT_12_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_12_MPORT_12_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_12_MPORT_12_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_12_MPORT_12_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_12_MPORT_140_en_pipe_0;
  reg [9:0] tensorFile_12_MPORT_140_addr_pipe_0;
  reg [63:0] tensorFile_13 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_13_MPORT_141_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_13_MPORT_141_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_13_MPORT_13_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_13_MPORT_13_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_13_MPORT_13_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_13_MPORT_13_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_13_MPORT_141_en_pipe_0;
  reg [9:0] tensorFile_13_MPORT_141_addr_pipe_0;
  reg [63:0] tensorFile_14 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_14_MPORT_142_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_14_MPORT_142_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_14_MPORT_14_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_14_MPORT_14_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_14_MPORT_14_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_14_MPORT_14_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_14_MPORT_142_en_pipe_0;
  reg [9:0] tensorFile_14_MPORT_142_addr_pipe_0;
  reg [63:0] tensorFile_15 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_15_MPORT_143_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_15_MPORT_143_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_15_MPORT_15_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_15_MPORT_15_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_15_MPORT_15_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_15_MPORT_15_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_15_MPORT_143_en_pipe_0;
  reg [9:0] tensorFile_15_MPORT_143_addr_pipe_0;
  reg [63:0] tensorFile_16 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_16_MPORT_144_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_16_MPORT_144_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_16_MPORT_16_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_16_MPORT_16_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_16_MPORT_16_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_16_MPORT_16_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_16_MPORT_144_en_pipe_0;
  reg [9:0] tensorFile_16_MPORT_144_addr_pipe_0;
  reg [63:0] tensorFile_17 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_17_MPORT_145_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_17_MPORT_145_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_17_MPORT_17_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_17_MPORT_17_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_17_MPORT_17_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_17_MPORT_17_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_17_MPORT_145_en_pipe_0;
  reg [9:0] tensorFile_17_MPORT_145_addr_pipe_0;
  reg [63:0] tensorFile_18 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_18_MPORT_146_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_18_MPORT_146_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_18_MPORT_18_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_18_MPORT_18_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_18_MPORT_18_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_18_MPORT_18_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_18_MPORT_146_en_pipe_0;
  reg [9:0] tensorFile_18_MPORT_146_addr_pipe_0;
  reg [63:0] tensorFile_19 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_19_MPORT_147_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_19_MPORT_147_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_19_MPORT_19_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_19_MPORT_19_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_19_MPORT_19_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_19_MPORT_19_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_19_MPORT_147_en_pipe_0;
  reg [9:0] tensorFile_19_MPORT_147_addr_pipe_0;
  reg [63:0] tensorFile_20 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_20_MPORT_148_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_20_MPORT_148_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_20_MPORT_20_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_20_MPORT_20_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_20_MPORT_20_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_20_MPORT_20_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_20_MPORT_148_en_pipe_0;
  reg [9:0] tensorFile_20_MPORT_148_addr_pipe_0;
  reg [63:0] tensorFile_21 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_21_MPORT_149_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_21_MPORT_149_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_21_MPORT_21_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_21_MPORT_21_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_21_MPORT_21_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_21_MPORT_21_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_21_MPORT_149_en_pipe_0;
  reg [9:0] tensorFile_21_MPORT_149_addr_pipe_0;
  reg [63:0] tensorFile_22 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_22_MPORT_150_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_22_MPORT_150_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_22_MPORT_22_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_22_MPORT_22_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_22_MPORT_22_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_22_MPORT_22_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_22_MPORT_150_en_pipe_0;
  reg [9:0] tensorFile_22_MPORT_150_addr_pipe_0;
  reg [63:0] tensorFile_23 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_23_MPORT_151_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_23_MPORT_151_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_23_MPORT_23_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_23_MPORT_23_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_23_MPORT_23_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_23_MPORT_23_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_23_MPORT_151_en_pipe_0;
  reg [9:0] tensorFile_23_MPORT_151_addr_pipe_0;
  reg [63:0] tensorFile_24 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_24_MPORT_152_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_24_MPORT_152_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_24_MPORT_24_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_24_MPORT_24_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_24_MPORT_24_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_24_MPORT_24_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_24_MPORT_152_en_pipe_0;
  reg [9:0] tensorFile_24_MPORT_152_addr_pipe_0;
  reg [63:0] tensorFile_25 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_25_MPORT_153_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_25_MPORT_153_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_25_MPORT_25_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_25_MPORT_25_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_25_MPORT_25_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_25_MPORT_25_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_25_MPORT_153_en_pipe_0;
  reg [9:0] tensorFile_25_MPORT_153_addr_pipe_0;
  reg [63:0] tensorFile_26 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_26_MPORT_154_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_26_MPORT_154_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_26_MPORT_26_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_26_MPORT_26_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_26_MPORT_26_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_26_MPORT_26_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_26_MPORT_154_en_pipe_0;
  reg [9:0] tensorFile_26_MPORT_154_addr_pipe_0;
  reg [63:0] tensorFile_27 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_27_MPORT_155_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_27_MPORT_155_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_27_MPORT_27_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_27_MPORT_27_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_27_MPORT_27_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_27_MPORT_27_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_27_MPORT_155_en_pipe_0;
  reg [9:0] tensorFile_27_MPORT_155_addr_pipe_0;
  reg [63:0] tensorFile_28 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_28_MPORT_156_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_28_MPORT_156_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_28_MPORT_28_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_28_MPORT_28_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_28_MPORT_28_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_28_MPORT_28_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_28_MPORT_156_en_pipe_0;
  reg [9:0] tensorFile_28_MPORT_156_addr_pipe_0;
  reg [63:0] tensorFile_29 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_29_MPORT_157_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_29_MPORT_157_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_29_MPORT_29_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_29_MPORT_29_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_29_MPORT_29_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_29_MPORT_29_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_29_MPORT_157_en_pipe_0;
  reg [9:0] tensorFile_29_MPORT_157_addr_pipe_0;
  reg [63:0] tensorFile_30 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_30_MPORT_158_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_30_MPORT_158_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_30_MPORT_30_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_30_MPORT_30_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_30_MPORT_30_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_30_MPORT_30_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_30_MPORT_158_en_pipe_0;
  reg [9:0] tensorFile_30_MPORT_158_addr_pipe_0;
  reg [63:0] tensorFile_31 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_31_MPORT_159_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_31_MPORT_159_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_31_MPORT_31_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_31_MPORT_31_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_31_MPORT_31_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_31_MPORT_31_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_31_MPORT_159_en_pipe_0;
  reg [9:0] tensorFile_31_MPORT_159_addr_pipe_0;
  reg [63:0] tensorFile_32 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_32_MPORT_160_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_32_MPORT_160_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_32_MPORT_32_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_32_MPORT_32_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_32_MPORT_32_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_32_MPORT_32_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_32_MPORT_160_en_pipe_0;
  reg [9:0] tensorFile_32_MPORT_160_addr_pipe_0;
  reg [63:0] tensorFile_33 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_33_MPORT_161_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_33_MPORT_161_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_33_MPORT_33_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_33_MPORT_33_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_33_MPORT_33_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_33_MPORT_33_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_33_MPORT_161_en_pipe_0;
  reg [9:0] tensorFile_33_MPORT_161_addr_pipe_0;
  reg [63:0] tensorFile_34 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_34_MPORT_162_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_34_MPORT_162_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_34_MPORT_34_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_34_MPORT_34_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_34_MPORT_34_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_34_MPORT_34_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_34_MPORT_162_en_pipe_0;
  reg [9:0] tensorFile_34_MPORT_162_addr_pipe_0;
  reg [63:0] tensorFile_35 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_35_MPORT_163_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_35_MPORT_163_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_35_MPORT_35_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_35_MPORT_35_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_35_MPORT_35_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_35_MPORT_35_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_35_MPORT_163_en_pipe_0;
  reg [9:0] tensorFile_35_MPORT_163_addr_pipe_0;
  reg [63:0] tensorFile_36 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_36_MPORT_164_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_36_MPORT_164_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_36_MPORT_36_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_36_MPORT_36_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_36_MPORT_36_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_36_MPORT_36_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_36_MPORT_164_en_pipe_0;
  reg [9:0] tensorFile_36_MPORT_164_addr_pipe_0;
  reg [63:0] tensorFile_37 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_37_MPORT_165_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_37_MPORT_165_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_37_MPORT_37_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_37_MPORT_37_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_37_MPORT_37_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_37_MPORT_37_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_37_MPORT_165_en_pipe_0;
  reg [9:0] tensorFile_37_MPORT_165_addr_pipe_0;
  reg [63:0] tensorFile_38 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_38_MPORT_166_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_38_MPORT_166_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_38_MPORT_38_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_38_MPORT_38_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_38_MPORT_38_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_38_MPORT_38_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_38_MPORT_166_en_pipe_0;
  reg [9:0] tensorFile_38_MPORT_166_addr_pipe_0;
  reg [63:0] tensorFile_39 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_39_MPORT_167_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_39_MPORT_167_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_39_MPORT_39_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_39_MPORT_39_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_39_MPORT_39_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_39_MPORT_39_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_39_MPORT_167_en_pipe_0;
  reg [9:0] tensorFile_39_MPORT_167_addr_pipe_0;
  reg [63:0] tensorFile_40 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_40_MPORT_168_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_40_MPORT_168_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_40_MPORT_40_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_40_MPORT_40_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_40_MPORT_40_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_40_MPORT_40_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_40_MPORT_168_en_pipe_0;
  reg [9:0] tensorFile_40_MPORT_168_addr_pipe_0;
  reg [63:0] tensorFile_41 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_41_MPORT_169_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_41_MPORT_169_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_41_MPORT_41_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_41_MPORT_41_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_41_MPORT_41_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_41_MPORT_41_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_41_MPORT_169_en_pipe_0;
  reg [9:0] tensorFile_41_MPORT_169_addr_pipe_0;
  reg [63:0] tensorFile_42 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_42_MPORT_170_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_42_MPORT_170_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_42_MPORT_42_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_42_MPORT_42_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_42_MPORT_42_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_42_MPORT_42_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_42_MPORT_170_en_pipe_0;
  reg [9:0] tensorFile_42_MPORT_170_addr_pipe_0;
  reg [63:0] tensorFile_43 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_43_MPORT_171_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_43_MPORT_171_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_43_MPORT_43_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_43_MPORT_43_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_43_MPORT_43_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_43_MPORT_43_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_43_MPORT_171_en_pipe_0;
  reg [9:0] tensorFile_43_MPORT_171_addr_pipe_0;
  reg [63:0] tensorFile_44 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_44_MPORT_172_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_44_MPORT_172_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_44_MPORT_44_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_44_MPORT_44_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_44_MPORT_44_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_44_MPORT_44_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_44_MPORT_172_en_pipe_0;
  reg [9:0] tensorFile_44_MPORT_172_addr_pipe_0;
  reg [63:0] tensorFile_45 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_45_MPORT_173_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_45_MPORT_173_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_45_MPORT_45_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_45_MPORT_45_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_45_MPORT_45_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_45_MPORT_45_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_45_MPORT_173_en_pipe_0;
  reg [9:0] tensorFile_45_MPORT_173_addr_pipe_0;
  reg [63:0] tensorFile_46 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_46_MPORT_174_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_46_MPORT_174_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_46_MPORT_46_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_46_MPORT_46_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_46_MPORT_46_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_46_MPORT_46_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_46_MPORT_174_en_pipe_0;
  reg [9:0] tensorFile_46_MPORT_174_addr_pipe_0;
  reg [63:0] tensorFile_47 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_47_MPORT_175_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_47_MPORT_175_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_47_MPORT_47_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_47_MPORT_47_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_47_MPORT_47_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_47_MPORT_47_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_47_MPORT_175_en_pipe_0;
  reg [9:0] tensorFile_47_MPORT_175_addr_pipe_0;
  reg [63:0] tensorFile_48 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_48_MPORT_176_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_48_MPORT_176_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_48_MPORT_48_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_48_MPORT_48_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_48_MPORT_48_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_48_MPORT_48_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_48_MPORT_176_en_pipe_0;
  reg [9:0] tensorFile_48_MPORT_176_addr_pipe_0;
  reg [63:0] tensorFile_49 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_49_MPORT_177_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_49_MPORT_177_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_49_MPORT_49_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_49_MPORT_49_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_49_MPORT_49_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_49_MPORT_49_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_49_MPORT_177_en_pipe_0;
  reg [9:0] tensorFile_49_MPORT_177_addr_pipe_0;
  reg [63:0] tensorFile_50 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_50_MPORT_178_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_50_MPORT_178_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_50_MPORT_50_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_50_MPORT_50_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_50_MPORT_50_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_50_MPORT_50_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_50_MPORT_178_en_pipe_0;
  reg [9:0] tensorFile_50_MPORT_178_addr_pipe_0;
  reg [63:0] tensorFile_51 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_51_MPORT_179_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_51_MPORT_179_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_51_MPORT_51_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_51_MPORT_51_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_51_MPORT_51_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_51_MPORT_51_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_51_MPORT_179_en_pipe_0;
  reg [9:0] tensorFile_51_MPORT_179_addr_pipe_0;
  reg [63:0] tensorFile_52 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_52_MPORT_180_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_52_MPORT_180_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_52_MPORT_52_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_52_MPORT_52_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_52_MPORT_52_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_52_MPORT_52_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_52_MPORT_180_en_pipe_0;
  reg [9:0] tensorFile_52_MPORT_180_addr_pipe_0;
  reg [63:0] tensorFile_53 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_53_MPORT_181_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_53_MPORT_181_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_53_MPORT_53_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_53_MPORT_53_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_53_MPORT_53_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_53_MPORT_53_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_53_MPORT_181_en_pipe_0;
  reg [9:0] tensorFile_53_MPORT_181_addr_pipe_0;
  reg [63:0] tensorFile_54 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_54_MPORT_182_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_54_MPORT_182_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_54_MPORT_54_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_54_MPORT_54_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_54_MPORT_54_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_54_MPORT_54_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_54_MPORT_182_en_pipe_0;
  reg [9:0] tensorFile_54_MPORT_182_addr_pipe_0;
  reg [63:0] tensorFile_55 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_55_MPORT_183_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_55_MPORT_183_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_55_MPORT_55_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_55_MPORT_55_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_55_MPORT_55_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_55_MPORT_55_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_55_MPORT_183_en_pipe_0;
  reg [9:0] tensorFile_55_MPORT_183_addr_pipe_0;
  reg [63:0] tensorFile_56 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_56_MPORT_184_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_56_MPORT_184_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_56_MPORT_56_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_56_MPORT_56_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_56_MPORT_56_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_56_MPORT_56_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_56_MPORT_184_en_pipe_0;
  reg [9:0] tensorFile_56_MPORT_184_addr_pipe_0;
  reg [63:0] tensorFile_57 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_57_MPORT_185_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_57_MPORT_185_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_57_MPORT_57_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_57_MPORT_57_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_57_MPORT_57_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_57_MPORT_57_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_57_MPORT_185_en_pipe_0;
  reg [9:0] tensorFile_57_MPORT_185_addr_pipe_0;
  reg [63:0] tensorFile_58 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_58_MPORT_186_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_58_MPORT_186_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_58_MPORT_58_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_58_MPORT_58_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_58_MPORT_58_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_58_MPORT_58_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_58_MPORT_186_en_pipe_0;
  reg [9:0] tensorFile_58_MPORT_186_addr_pipe_0;
  reg [63:0] tensorFile_59 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_59_MPORT_187_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_59_MPORT_187_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_59_MPORT_59_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_59_MPORT_59_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_59_MPORT_59_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_59_MPORT_59_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_59_MPORT_187_en_pipe_0;
  reg [9:0] tensorFile_59_MPORT_187_addr_pipe_0;
  reg [63:0] tensorFile_60 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_60_MPORT_188_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_60_MPORT_188_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_60_MPORT_60_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_60_MPORT_60_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_60_MPORT_60_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_60_MPORT_60_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_60_MPORT_188_en_pipe_0;
  reg [9:0] tensorFile_60_MPORT_188_addr_pipe_0;
  reg [63:0] tensorFile_61 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_61_MPORT_189_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_61_MPORT_189_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_61_MPORT_61_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_61_MPORT_61_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_61_MPORT_61_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_61_MPORT_61_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_61_MPORT_189_en_pipe_0;
  reg [9:0] tensorFile_61_MPORT_189_addr_pipe_0;
  reg [63:0] tensorFile_62 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_62_MPORT_190_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_62_MPORT_190_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_62_MPORT_62_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_62_MPORT_62_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_62_MPORT_62_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_62_MPORT_62_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_62_MPORT_190_en_pipe_0;
  reg [9:0] tensorFile_62_MPORT_190_addr_pipe_0;
  reg [63:0] tensorFile_63 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_63_MPORT_191_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_63_MPORT_191_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_63_MPORT_63_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_63_MPORT_63_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_63_MPORT_63_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_63_MPORT_63_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_63_MPORT_191_en_pipe_0;
  reg [9:0] tensorFile_63_MPORT_191_addr_pipe_0;
  reg [63:0] tensorFile_64 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_64_MPORT_192_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_64_MPORT_192_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_64_MPORT_64_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_64_MPORT_64_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_64_MPORT_64_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_64_MPORT_64_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_64_MPORT_192_en_pipe_0;
  reg [9:0] tensorFile_64_MPORT_192_addr_pipe_0;
  reg [63:0] tensorFile_65 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_65_MPORT_193_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_65_MPORT_193_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_65_MPORT_65_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_65_MPORT_65_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_65_MPORT_65_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_65_MPORT_65_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_65_MPORT_193_en_pipe_0;
  reg [9:0] tensorFile_65_MPORT_193_addr_pipe_0;
  reg [63:0] tensorFile_66 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_66_MPORT_194_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_66_MPORT_194_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_66_MPORT_66_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_66_MPORT_66_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_66_MPORT_66_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_66_MPORT_66_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_66_MPORT_194_en_pipe_0;
  reg [9:0] tensorFile_66_MPORT_194_addr_pipe_0;
  reg [63:0] tensorFile_67 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_67_MPORT_195_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_67_MPORT_195_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_67_MPORT_67_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_67_MPORT_67_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_67_MPORT_67_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_67_MPORT_67_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_67_MPORT_195_en_pipe_0;
  reg [9:0] tensorFile_67_MPORT_195_addr_pipe_0;
  reg [63:0] tensorFile_68 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_68_MPORT_196_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_68_MPORT_196_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_68_MPORT_68_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_68_MPORT_68_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_68_MPORT_68_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_68_MPORT_68_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_68_MPORT_196_en_pipe_0;
  reg [9:0] tensorFile_68_MPORT_196_addr_pipe_0;
  reg [63:0] tensorFile_69 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_69_MPORT_197_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_69_MPORT_197_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_69_MPORT_69_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_69_MPORT_69_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_69_MPORT_69_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_69_MPORT_69_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_69_MPORT_197_en_pipe_0;
  reg [9:0] tensorFile_69_MPORT_197_addr_pipe_0;
  reg [63:0] tensorFile_70 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_70_MPORT_198_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_70_MPORT_198_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_70_MPORT_70_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_70_MPORT_70_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_70_MPORT_70_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_70_MPORT_70_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_70_MPORT_198_en_pipe_0;
  reg [9:0] tensorFile_70_MPORT_198_addr_pipe_0;
  reg [63:0] tensorFile_71 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_71_MPORT_199_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_71_MPORT_199_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_71_MPORT_71_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_71_MPORT_71_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_71_MPORT_71_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_71_MPORT_71_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_71_MPORT_199_en_pipe_0;
  reg [9:0] tensorFile_71_MPORT_199_addr_pipe_0;
  reg [63:0] tensorFile_72 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_72_MPORT_200_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_72_MPORT_200_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_72_MPORT_72_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_72_MPORT_72_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_72_MPORT_72_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_72_MPORT_72_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_72_MPORT_200_en_pipe_0;
  reg [9:0] tensorFile_72_MPORT_200_addr_pipe_0;
  reg [63:0] tensorFile_73 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_73_MPORT_201_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_73_MPORT_201_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_73_MPORT_73_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_73_MPORT_73_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_73_MPORT_73_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_73_MPORT_73_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_73_MPORT_201_en_pipe_0;
  reg [9:0] tensorFile_73_MPORT_201_addr_pipe_0;
  reg [63:0] tensorFile_74 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_74_MPORT_202_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_74_MPORT_202_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_74_MPORT_74_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_74_MPORT_74_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_74_MPORT_74_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_74_MPORT_74_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_74_MPORT_202_en_pipe_0;
  reg [9:0] tensorFile_74_MPORT_202_addr_pipe_0;
  reg [63:0] tensorFile_75 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_75_MPORT_203_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_75_MPORT_203_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_75_MPORT_75_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_75_MPORT_75_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_75_MPORT_75_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_75_MPORT_75_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_75_MPORT_203_en_pipe_0;
  reg [9:0] tensorFile_75_MPORT_203_addr_pipe_0;
  reg [63:0] tensorFile_76 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_76_MPORT_204_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_76_MPORT_204_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_76_MPORT_76_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_76_MPORT_76_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_76_MPORT_76_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_76_MPORT_76_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_76_MPORT_204_en_pipe_0;
  reg [9:0] tensorFile_76_MPORT_204_addr_pipe_0;
  reg [63:0] tensorFile_77 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_77_MPORT_205_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_77_MPORT_205_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_77_MPORT_77_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_77_MPORT_77_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_77_MPORT_77_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_77_MPORT_77_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_77_MPORT_205_en_pipe_0;
  reg [9:0] tensorFile_77_MPORT_205_addr_pipe_0;
  reg [63:0] tensorFile_78 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_78_MPORT_206_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_78_MPORT_206_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_78_MPORT_78_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_78_MPORT_78_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_78_MPORT_78_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_78_MPORT_78_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_78_MPORT_206_en_pipe_0;
  reg [9:0] tensorFile_78_MPORT_206_addr_pipe_0;
  reg [63:0] tensorFile_79 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_79_MPORT_207_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_79_MPORT_207_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_79_MPORT_79_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_79_MPORT_79_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_79_MPORT_79_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_79_MPORT_79_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_79_MPORT_207_en_pipe_0;
  reg [9:0] tensorFile_79_MPORT_207_addr_pipe_0;
  reg [63:0] tensorFile_80 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_80_MPORT_208_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_80_MPORT_208_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_80_MPORT_80_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_80_MPORT_80_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_80_MPORT_80_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_80_MPORT_80_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_80_MPORT_208_en_pipe_0;
  reg [9:0] tensorFile_80_MPORT_208_addr_pipe_0;
  reg [63:0] tensorFile_81 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_81_MPORT_209_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_81_MPORT_209_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_81_MPORT_81_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_81_MPORT_81_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_81_MPORT_81_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_81_MPORT_81_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_81_MPORT_209_en_pipe_0;
  reg [9:0] tensorFile_81_MPORT_209_addr_pipe_0;
  reg [63:0] tensorFile_82 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_82_MPORT_210_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_82_MPORT_210_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_82_MPORT_82_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_82_MPORT_82_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_82_MPORT_82_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_82_MPORT_82_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_82_MPORT_210_en_pipe_0;
  reg [9:0] tensorFile_82_MPORT_210_addr_pipe_0;
  reg [63:0] tensorFile_83 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_83_MPORT_211_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_83_MPORT_211_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_83_MPORT_83_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_83_MPORT_83_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_83_MPORT_83_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_83_MPORT_83_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_83_MPORT_211_en_pipe_0;
  reg [9:0] tensorFile_83_MPORT_211_addr_pipe_0;
  reg [63:0] tensorFile_84 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_84_MPORT_212_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_84_MPORT_212_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_84_MPORT_84_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_84_MPORT_84_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_84_MPORT_84_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_84_MPORT_84_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_84_MPORT_212_en_pipe_0;
  reg [9:0] tensorFile_84_MPORT_212_addr_pipe_0;
  reg [63:0] tensorFile_85 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_85_MPORT_213_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_85_MPORT_213_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_85_MPORT_85_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_85_MPORT_85_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_85_MPORT_85_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_85_MPORT_85_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_85_MPORT_213_en_pipe_0;
  reg [9:0] tensorFile_85_MPORT_213_addr_pipe_0;
  reg [63:0] tensorFile_86 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_86_MPORT_214_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_86_MPORT_214_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_86_MPORT_86_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_86_MPORT_86_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_86_MPORT_86_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_86_MPORT_86_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_86_MPORT_214_en_pipe_0;
  reg [9:0] tensorFile_86_MPORT_214_addr_pipe_0;
  reg [63:0] tensorFile_87 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_87_MPORT_215_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_87_MPORT_215_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_87_MPORT_87_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_87_MPORT_87_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_87_MPORT_87_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_87_MPORT_87_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_87_MPORT_215_en_pipe_0;
  reg [9:0] tensorFile_87_MPORT_215_addr_pipe_0;
  reg [63:0] tensorFile_88 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_88_MPORT_216_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_88_MPORT_216_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_88_MPORT_88_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_88_MPORT_88_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_88_MPORT_88_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_88_MPORT_88_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_88_MPORT_216_en_pipe_0;
  reg [9:0] tensorFile_88_MPORT_216_addr_pipe_0;
  reg [63:0] tensorFile_89 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_89_MPORT_217_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_89_MPORT_217_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_89_MPORT_89_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_89_MPORT_89_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_89_MPORT_89_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_89_MPORT_89_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_89_MPORT_217_en_pipe_0;
  reg [9:0] tensorFile_89_MPORT_217_addr_pipe_0;
  reg [63:0] tensorFile_90 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_90_MPORT_218_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_90_MPORT_218_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_90_MPORT_90_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_90_MPORT_90_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_90_MPORT_90_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_90_MPORT_90_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_90_MPORT_218_en_pipe_0;
  reg [9:0] tensorFile_90_MPORT_218_addr_pipe_0;
  reg [63:0] tensorFile_91 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_91_MPORT_219_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_91_MPORT_219_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_91_MPORT_91_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_91_MPORT_91_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_91_MPORT_91_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_91_MPORT_91_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_91_MPORT_219_en_pipe_0;
  reg [9:0] tensorFile_91_MPORT_219_addr_pipe_0;
  reg [63:0] tensorFile_92 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_92_MPORT_220_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_92_MPORT_220_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_92_MPORT_92_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_92_MPORT_92_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_92_MPORT_92_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_92_MPORT_92_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_92_MPORT_220_en_pipe_0;
  reg [9:0] tensorFile_92_MPORT_220_addr_pipe_0;
  reg [63:0] tensorFile_93 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_93_MPORT_221_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_93_MPORT_221_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_93_MPORT_93_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_93_MPORT_93_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_93_MPORT_93_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_93_MPORT_93_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_93_MPORT_221_en_pipe_0;
  reg [9:0] tensorFile_93_MPORT_221_addr_pipe_0;
  reg [63:0] tensorFile_94 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_94_MPORT_222_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_94_MPORT_222_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_94_MPORT_94_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_94_MPORT_94_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_94_MPORT_94_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_94_MPORT_94_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_94_MPORT_222_en_pipe_0;
  reg [9:0] tensorFile_94_MPORT_222_addr_pipe_0;
  reg [63:0] tensorFile_95 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_95_MPORT_223_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_95_MPORT_223_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_95_MPORT_95_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_95_MPORT_95_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_95_MPORT_95_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_95_MPORT_95_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_95_MPORT_223_en_pipe_0;
  reg [9:0] tensorFile_95_MPORT_223_addr_pipe_0;
  reg [63:0] tensorFile_96 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_96_MPORT_224_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_96_MPORT_224_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_96_MPORT_96_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_96_MPORT_96_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_96_MPORT_96_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_96_MPORT_96_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_96_MPORT_224_en_pipe_0;
  reg [9:0] tensorFile_96_MPORT_224_addr_pipe_0;
  reg [63:0] tensorFile_97 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_97_MPORT_225_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_97_MPORT_225_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_97_MPORT_97_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_97_MPORT_97_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_97_MPORT_97_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_97_MPORT_97_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_97_MPORT_225_en_pipe_0;
  reg [9:0] tensorFile_97_MPORT_225_addr_pipe_0;
  reg [63:0] tensorFile_98 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_98_MPORT_226_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_98_MPORT_226_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_98_MPORT_98_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_98_MPORT_98_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_98_MPORT_98_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_98_MPORT_98_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_98_MPORT_226_en_pipe_0;
  reg [9:0] tensorFile_98_MPORT_226_addr_pipe_0;
  reg [63:0] tensorFile_99 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_99_MPORT_227_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_99_MPORT_227_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_99_MPORT_99_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_99_MPORT_99_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_99_MPORT_99_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_99_MPORT_99_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_99_MPORT_227_en_pipe_0;
  reg [9:0] tensorFile_99_MPORT_227_addr_pipe_0;
  reg [63:0] tensorFile_100 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_100_MPORT_228_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_100_MPORT_228_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_100_MPORT_100_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_100_MPORT_100_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_100_MPORT_100_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_100_MPORT_100_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_100_MPORT_228_en_pipe_0;
  reg [9:0] tensorFile_100_MPORT_228_addr_pipe_0;
  reg [63:0] tensorFile_101 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_101_MPORT_229_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_101_MPORT_229_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_101_MPORT_101_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_101_MPORT_101_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_101_MPORT_101_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_101_MPORT_101_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_101_MPORT_229_en_pipe_0;
  reg [9:0] tensorFile_101_MPORT_229_addr_pipe_0;
  reg [63:0] tensorFile_102 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_102_MPORT_230_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_102_MPORT_230_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_102_MPORT_102_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_102_MPORT_102_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_102_MPORT_102_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_102_MPORT_102_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_102_MPORT_230_en_pipe_0;
  reg [9:0] tensorFile_102_MPORT_230_addr_pipe_0;
  reg [63:0] tensorFile_103 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_103_MPORT_231_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_103_MPORT_231_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_103_MPORT_103_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_103_MPORT_103_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_103_MPORT_103_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_103_MPORT_103_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_103_MPORT_231_en_pipe_0;
  reg [9:0] tensorFile_103_MPORT_231_addr_pipe_0;
  reg [63:0] tensorFile_104 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_104_MPORT_232_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_104_MPORT_232_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_104_MPORT_104_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_104_MPORT_104_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_104_MPORT_104_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_104_MPORT_104_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_104_MPORT_232_en_pipe_0;
  reg [9:0] tensorFile_104_MPORT_232_addr_pipe_0;
  reg [63:0] tensorFile_105 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_105_MPORT_233_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_105_MPORT_233_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_105_MPORT_105_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_105_MPORT_105_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_105_MPORT_105_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_105_MPORT_105_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_105_MPORT_233_en_pipe_0;
  reg [9:0] tensorFile_105_MPORT_233_addr_pipe_0;
  reg [63:0] tensorFile_106 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_106_MPORT_234_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_106_MPORT_234_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_106_MPORT_106_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_106_MPORT_106_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_106_MPORT_106_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_106_MPORT_106_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_106_MPORT_234_en_pipe_0;
  reg [9:0] tensorFile_106_MPORT_234_addr_pipe_0;
  reg [63:0] tensorFile_107 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_107_MPORT_235_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_107_MPORT_235_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_107_MPORT_107_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_107_MPORT_107_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_107_MPORT_107_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_107_MPORT_107_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_107_MPORT_235_en_pipe_0;
  reg [9:0] tensorFile_107_MPORT_235_addr_pipe_0;
  reg [63:0] tensorFile_108 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_108_MPORT_236_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_108_MPORT_236_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_108_MPORT_108_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_108_MPORT_108_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_108_MPORT_108_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_108_MPORT_108_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_108_MPORT_236_en_pipe_0;
  reg [9:0] tensorFile_108_MPORT_236_addr_pipe_0;
  reg [63:0] tensorFile_109 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_109_MPORT_237_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_109_MPORT_237_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_109_MPORT_109_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_109_MPORT_109_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_109_MPORT_109_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_109_MPORT_109_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_109_MPORT_237_en_pipe_0;
  reg [9:0] tensorFile_109_MPORT_237_addr_pipe_0;
  reg [63:0] tensorFile_110 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_110_MPORT_238_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_110_MPORT_238_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_110_MPORT_110_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_110_MPORT_110_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_110_MPORT_110_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_110_MPORT_110_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_110_MPORT_238_en_pipe_0;
  reg [9:0] tensorFile_110_MPORT_238_addr_pipe_0;
  reg [63:0] tensorFile_111 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_111_MPORT_239_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_111_MPORT_239_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_111_MPORT_111_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_111_MPORT_111_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_111_MPORT_111_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_111_MPORT_111_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_111_MPORT_239_en_pipe_0;
  reg [9:0] tensorFile_111_MPORT_239_addr_pipe_0;
  reg [63:0] tensorFile_112 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_112_MPORT_240_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_112_MPORT_240_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_112_MPORT_112_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_112_MPORT_112_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_112_MPORT_112_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_112_MPORT_112_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_112_MPORT_240_en_pipe_0;
  reg [9:0] tensorFile_112_MPORT_240_addr_pipe_0;
  reg [63:0] tensorFile_113 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_113_MPORT_241_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_113_MPORT_241_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_113_MPORT_113_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_113_MPORT_113_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_113_MPORT_113_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_113_MPORT_113_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_113_MPORT_241_en_pipe_0;
  reg [9:0] tensorFile_113_MPORT_241_addr_pipe_0;
  reg [63:0] tensorFile_114 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_114_MPORT_242_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_114_MPORT_242_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_114_MPORT_114_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_114_MPORT_114_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_114_MPORT_114_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_114_MPORT_114_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_114_MPORT_242_en_pipe_0;
  reg [9:0] tensorFile_114_MPORT_242_addr_pipe_0;
  reg [63:0] tensorFile_115 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_115_MPORT_243_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_115_MPORT_243_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_115_MPORT_115_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_115_MPORT_115_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_115_MPORT_115_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_115_MPORT_115_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_115_MPORT_243_en_pipe_0;
  reg [9:0] tensorFile_115_MPORT_243_addr_pipe_0;
  reg [63:0] tensorFile_116 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_116_MPORT_244_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_116_MPORT_244_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_116_MPORT_116_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_116_MPORT_116_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_116_MPORT_116_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_116_MPORT_116_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_116_MPORT_244_en_pipe_0;
  reg [9:0] tensorFile_116_MPORT_244_addr_pipe_0;
  reg [63:0] tensorFile_117 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_117_MPORT_245_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_117_MPORT_245_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_117_MPORT_117_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_117_MPORT_117_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_117_MPORT_117_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_117_MPORT_117_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_117_MPORT_245_en_pipe_0;
  reg [9:0] tensorFile_117_MPORT_245_addr_pipe_0;
  reg [63:0] tensorFile_118 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_118_MPORT_246_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_118_MPORT_246_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_118_MPORT_118_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_118_MPORT_118_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_118_MPORT_118_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_118_MPORT_118_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_118_MPORT_246_en_pipe_0;
  reg [9:0] tensorFile_118_MPORT_246_addr_pipe_0;
  reg [63:0] tensorFile_119 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_119_MPORT_247_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_119_MPORT_247_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_119_MPORT_119_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_119_MPORT_119_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_119_MPORT_119_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_119_MPORT_119_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_119_MPORT_247_en_pipe_0;
  reg [9:0] tensorFile_119_MPORT_247_addr_pipe_0;
  reg [63:0] tensorFile_120 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_120_MPORT_248_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_120_MPORT_248_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_120_MPORT_120_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_120_MPORT_120_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_120_MPORT_120_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_120_MPORT_120_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_120_MPORT_248_en_pipe_0;
  reg [9:0] tensorFile_120_MPORT_248_addr_pipe_0;
  reg [63:0] tensorFile_121 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_121_MPORT_249_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_121_MPORT_249_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_121_MPORT_121_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_121_MPORT_121_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_121_MPORT_121_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_121_MPORT_121_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_121_MPORT_249_en_pipe_0;
  reg [9:0] tensorFile_121_MPORT_249_addr_pipe_0;
  reg [63:0] tensorFile_122 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_122_MPORT_250_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_122_MPORT_250_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_122_MPORT_122_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_122_MPORT_122_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_122_MPORT_122_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_122_MPORT_122_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_122_MPORT_250_en_pipe_0;
  reg [9:0] tensorFile_122_MPORT_250_addr_pipe_0;
  reg [63:0] tensorFile_123 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_123_MPORT_251_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_123_MPORT_251_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_123_MPORT_123_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_123_MPORT_123_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_123_MPORT_123_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_123_MPORT_123_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_123_MPORT_251_en_pipe_0;
  reg [9:0] tensorFile_123_MPORT_251_addr_pipe_0;
  reg [63:0] tensorFile_124 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_124_MPORT_252_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_124_MPORT_252_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_124_MPORT_124_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_124_MPORT_124_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_124_MPORT_124_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_124_MPORT_124_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_124_MPORT_252_en_pipe_0;
  reg [9:0] tensorFile_124_MPORT_252_addr_pipe_0;
  reg [63:0] tensorFile_125 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_125_MPORT_253_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_125_MPORT_253_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_125_MPORT_125_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_125_MPORT_125_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_125_MPORT_125_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_125_MPORT_125_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_125_MPORT_253_en_pipe_0;
  reg [9:0] tensorFile_125_MPORT_253_addr_pipe_0;
  reg [63:0] tensorFile_126 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_126_MPORT_254_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_126_MPORT_254_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_126_MPORT_126_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_126_MPORT_126_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_126_MPORT_126_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_126_MPORT_126_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_126_MPORT_254_en_pipe_0;
  reg [9:0] tensorFile_126_MPORT_254_addr_pipe_0;
  reg [63:0] tensorFile_127 [0:1023]; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_127_MPORT_255_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_127_MPORT_255_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_127_MPORT_127_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [9:0] tensorFile_127_MPORT_127_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_127_MPORT_127_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_127_MPORT_127_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_127_MPORT_255_en_pipe_0;
  reg [9:0] tensorFile_127_MPORT_255_addr_pipe_0;
  reg  state; // @[TensorLoadNarrowVME.scala 54:22]
  reg [16:0] blocksInFlight; // @[TensorLoadNarrowVME.scala 87:27]
  wire  loadDone = blocksInFlight == 17'h0 & vmeCmd_io_done & state; // @[TensorLoadNarrowVME.scala 292:57]
  wire  localDone = loadDone & fillPadding_io_done; // @[TensorLoadNarrowVME.scala 293:25]
  wire  _GEN_0 = localDone ? 1'h0 : state; // @[TensorLoadNarrowVME.scala 61:25 TensorLoadNarrowVME.scala 62:11 TensorLoadNarrowVME.scala 54:22]
  wire  _GEN_1 = io_start | _GEN_0; // @[TensorLoadNarrowVME.scala 59:18 TensorLoadNarrowVME.scala 60:11]
  reg [63:0] vmeDataBitsPipe_data; // @[TensorLoadNarrowVME.scala 67:32]
  reg [20:0] vmeDataBitsPipe_tag; // @[TensorLoadNarrowVME.scala 67:32]
  reg  vmeDataValidPipe; // @[TensorLoadNarrowVME.scala 68:33]
  reg  vmeDataReadyPipe; // @[TensorLoadNarrowVME.scala 69:33]
  wire  vmeDataFirePipe = vmeDataValidPipe & vmeDataReadyPipe; // @[TensorLoadNarrowVME.scala 70:42]
  wire  _T = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[Decoupled.scala 40:37]
  wire  _T_1 = state & _T; // @[TensorLoadNarrowVME.scala 90:21]
  wire  _T_3 = state & _T & ~vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 90:45]
  wire [16:0] _GEN_778 = {{8'd0}, vmeCmd_io_readLen}; // @[TensorLoadNarrowVME.scala 91:38]
  wire [16:0] _blocksInFlight_T_1 = blocksInFlight + _GEN_778; // @[TensorLoadNarrowVME.scala 91:38]
  wire  _T_6 = _T_1 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 92:45]
  wire [16:0] _blocksInFlight_T_5 = _blocksInFlight_T_1 - 17'h1; // @[TensorLoadNarrowVME.scala 93:48]
  wire  _T_10 = state & ~_T & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 94:46]
  wire [16:0] _blocksInFlight_T_7 = blocksInFlight - 17'h1; // @[TensorLoadNarrowVME.scala 96:38]
  reg [127:0] fillPadding_io_inst_REG; // @[TensorLoadNarrowVME.scala 121:33]
  reg  fillPadding_io_start_REG; // @[TensorLoadNarrowVME.scala 122:34]
  wire [9:0] waddrTensInstrTmp = fillPadding_io_tensorIdx_valid ? fillPadding_io_tensorIdx_bits : readData_io_idx; // @[TensorLoadNarrowVME.scala 166:30]
  wire  _waddr_0_T = ~state; // @[TensorLoadNarrowVME.scala 186:27]
  wire  wenTensInstr_0 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h0 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_1 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h1 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_2 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h2 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_3 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h3 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_4 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h4 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_5 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h5 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_6 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h6 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_7 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h7 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_8 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h8 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_9 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h9 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_10 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'ha & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_11 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'hb & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_12 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'hc & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_13 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'hd & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_14 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'he & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_15 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'hf & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_16 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h10 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_17 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h11 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_18 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h12 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_19 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h13 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_20 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h14 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_21 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h15 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_22 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h16 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_23 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h17 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_24 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h18 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_25 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h19 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_26 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h1a & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_27 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h1b & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_28 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h1c & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_29 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h1d & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_30 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h1e & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_31 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h1f & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_32 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h20 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_33 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h21 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_34 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h22 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_35 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h23 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_36 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h24 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_37 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h25 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_38 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h26 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_39 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h27 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_40 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h28 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_41 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h29 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_42 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h2a & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_43 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h2b & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_44 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h2c & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_45 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h2d & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_46 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h2e & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_47 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h2f & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_48 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h30 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_49 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h31 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_50 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h32 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_51 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h33 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_52 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h34 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_53 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h35 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_54 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h36 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_55 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h37 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_56 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h38 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_57 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h39 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_58 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h3a & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_59 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h3b & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_60 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h3c & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_61 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h3d & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_62 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h3e & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_63 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h3f & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_64 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h40 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_65 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h41 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_66 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h42 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_67 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h43 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_68 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h44 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_69 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h45 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_70 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h46 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_71 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h47 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_72 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h48 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_73 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h49 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_74 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h4a & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_75 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h4b & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_76 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h4c & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_77 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h4d & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_78 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h4e & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_79 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h4f & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_80 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h50 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_81 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h51 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_82 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h52 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_83 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h53 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_84 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h54 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_85 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h55 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_86 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h56 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_87 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h57 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_88 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h58 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_89 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h59 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_90 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h5a & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_91 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h5b & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_92 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h5c & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_93 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h5d & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_94 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h5e & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_95 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h5f & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_96 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h60 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_97 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h61 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_98 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h62 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_99 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h63 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_100 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h64 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_101 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h65 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_102 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h66 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_103 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h67 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_104 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h68 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_105 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h69 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_106 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h6a & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_107 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h6b & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_108 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h6c & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_109 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h6d & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_110 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h6e & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_111 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h6f & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_112 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h70 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_113 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h71 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_114 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h72 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_115 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h73 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_116 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h74 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_117 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h75 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_118 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h76 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_119 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h77 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_120 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h78 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_121 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h79 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_122 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h7a & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_123 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h7b & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_124 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h7c & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_125 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h7d & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_126 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h7e & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_127 = fillPadding_io_tensorIdx_valid | readData_io_col == 7'h7f & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire [63:0] wdataTensInstr_0 = fillPadding_io_tensorIdx_valid ? 64'h0 : vmeDataBitsPipe_data; // @[TensorLoadNarrowVME.scala 234:29]
  reg  rvalid; // @[Reg.scala 27:20]
  wire [63:0] _WIRE_128_1 = tensorFile_1_MPORT_129_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_0 = tensorFile_0_MPORT_128_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_3 = tensorFile_3_MPORT_131_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_2 = tensorFile_2_MPORT_130_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_5 = tensorFile_5_MPORT_133_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_4 = tensorFile_4_MPORT_132_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_7 = tensorFile_7_MPORT_135_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_6 = tensorFile_6_MPORT_134_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [511:0] lo_lo_lo_lo = {_WIRE_128_7,_WIRE_128_6,_WIRE_128_5,_WIRE_128_4,_WIRE_128_3,_WIRE_128_2,_WIRE_128_1,
    _WIRE_128_0}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_9 = tensorFile_9_MPORT_137_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_8 = tensorFile_8_MPORT_136_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_11 = tensorFile_11_MPORT_139_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_10 = tensorFile_10_MPORT_138_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_13 = tensorFile_13_MPORT_141_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_12 = tensorFile_12_MPORT_140_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_15 = tensorFile_15_MPORT_143_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_14 = tensorFile_14_MPORT_142_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [1023:0] lo_lo_lo = {_WIRE_128_15,_WIRE_128_14,_WIRE_128_13,_WIRE_128_12,_WIRE_128_11,_WIRE_128_10,_WIRE_128_9,
    _WIRE_128_8,lo_lo_lo_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_17 = tensorFile_17_MPORT_145_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_16 = tensorFile_16_MPORT_144_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_19 = tensorFile_19_MPORT_147_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_18 = tensorFile_18_MPORT_146_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_21 = tensorFile_21_MPORT_149_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_20 = tensorFile_20_MPORT_148_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_23 = tensorFile_23_MPORT_151_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_22 = tensorFile_22_MPORT_150_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [511:0] lo_lo_hi_lo = {_WIRE_128_23,_WIRE_128_22,_WIRE_128_21,_WIRE_128_20,_WIRE_128_19,_WIRE_128_18,_WIRE_128_17
    ,_WIRE_128_16}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_25 = tensorFile_25_MPORT_153_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_24 = tensorFile_24_MPORT_152_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_27 = tensorFile_27_MPORT_155_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_26 = tensorFile_26_MPORT_154_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_29 = tensorFile_29_MPORT_157_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_28 = tensorFile_28_MPORT_156_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_31 = tensorFile_31_MPORT_159_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_30 = tensorFile_30_MPORT_158_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [2047:0] lo_lo = {_WIRE_128_31,_WIRE_128_30,_WIRE_128_29,_WIRE_128_28,_WIRE_128_27,_WIRE_128_26,_WIRE_128_25,
    _WIRE_128_24,lo_lo_hi_lo,lo_lo_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_33 = tensorFile_33_MPORT_161_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_32 = tensorFile_32_MPORT_160_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_35 = tensorFile_35_MPORT_163_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_34 = tensorFile_34_MPORT_162_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_37 = tensorFile_37_MPORT_165_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_36 = tensorFile_36_MPORT_164_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_39 = tensorFile_39_MPORT_167_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_38 = tensorFile_38_MPORT_166_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [511:0] lo_hi_lo_lo = {_WIRE_128_39,_WIRE_128_38,_WIRE_128_37,_WIRE_128_36,_WIRE_128_35,_WIRE_128_34,_WIRE_128_33
    ,_WIRE_128_32}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_41 = tensorFile_41_MPORT_169_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_40 = tensorFile_40_MPORT_168_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_43 = tensorFile_43_MPORT_171_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_42 = tensorFile_42_MPORT_170_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_45 = tensorFile_45_MPORT_173_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_44 = tensorFile_44_MPORT_172_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_47 = tensorFile_47_MPORT_175_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_46 = tensorFile_46_MPORT_174_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [1023:0] lo_hi_lo = {_WIRE_128_47,_WIRE_128_46,_WIRE_128_45,_WIRE_128_44,_WIRE_128_43,_WIRE_128_42,_WIRE_128_41,
    _WIRE_128_40,lo_hi_lo_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_49 = tensorFile_49_MPORT_177_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_48 = tensorFile_48_MPORT_176_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_51 = tensorFile_51_MPORT_179_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_50 = tensorFile_50_MPORT_178_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_53 = tensorFile_53_MPORT_181_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_52 = tensorFile_52_MPORT_180_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_55 = tensorFile_55_MPORT_183_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_54 = tensorFile_54_MPORT_182_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [511:0] lo_hi_hi_lo = {_WIRE_128_55,_WIRE_128_54,_WIRE_128_53,_WIRE_128_52,_WIRE_128_51,_WIRE_128_50,_WIRE_128_49
    ,_WIRE_128_48}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_57 = tensorFile_57_MPORT_185_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_56 = tensorFile_56_MPORT_184_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_59 = tensorFile_59_MPORT_187_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_58 = tensorFile_58_MPORT_186_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_61 = tensorFile_61_MPORT_189_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_60 = tensorFile_60_MPORT_188_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_63 = tensorFile_63_MPORT_191_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_62 = tensorFile_62_MPORT_190_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [2047:0] lo_hi = {_WIRE_128_63,_WIRE_128_62,_WIRE_128_61,_WIRE_128_60,_WIRE_128_59,_WIRE_128_58,_WIRE_128_57,
    _WIRE_128_56,lo_hi_hi_lo,lo_hi_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_65 = tensorFile_65_MPORT_193_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_64 = tensorFile_64_MPORT_192_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_67 = tensorFile_67_MPORT_195_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_66 = tensorFile_66_MPORT_194_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_69 = tensorFile_69_MPORT_197_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_68 = tensorFile_68_MPORT_196_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_71 = tensorFile_71_MPORT_199_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_70 = tensorFile_70_MPORT_198_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [511:0] hi_lo_lo_lo = {_WIRE_128_71,_WIRE_128_70,_WIRE_128_69,_WIRE_128_68,_WIRE_128_67,_WIRE_128_66,_WIRE_128_65
    ,_WIRE_128_64}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_73 = tensorFile_73_MPORT_201_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_72 = tensorFile_72_MPORT_200_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_75 = tensorFile_75_MPORT_203_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_74 = tensorFile_74_MPORT_202_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_77 = tensorFile_77_MPORT_205_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_76 = tensorFile_76_MPORT_204_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_79 = tensorFile_79_MPORT_207_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_78 = tensorFile_78_MPORT_206_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [1023:0] hi_lo_lo = {_WIRE_128_79,_WIRE_128_78,_WIRE_128_77,_WIRE_128_76,_WIRE_128_75,_WIRE_128_74,_WIRE_128_73,
    _WIRE_128_72,hi_lo_lo_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_81 = tensorFile_81_MPORT_209_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_80 = tensorFile_80_MPORT_208_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_83 = tensorFile_83_MPORT_211_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_82 = tensorFile_82_MPORT_210_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_85 = tensorFile_85_MPORT_213_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_84 = tensorFile_84_MPORT_212_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_87 = tensorFile_87_MPORT_215_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_86 = tensorFile_86_MPORT_214_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [511:0] hi_lo_hi_lo = {_WIRE_128_87,_WIRE_128_86,_WIRE_128_85,_WIRE_128_84,_WIRE_128_83,_WIRE_128_82,_WIRE_128_81
    ,_WIRE_128_80}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_89 = tensorFile_89_MPORT_217_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_88 = tensorFile_88_MPORT_216_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_91 = tensorFile_91_MPORT_219_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_90 = tensorFile_90_MPORT_218_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_93 = tensorFile_93_MPORT_221_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_92 = tensorFile_92_MPORT_220_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_95 = tensorFile_95_MPORT_223_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_94 = tensorFile_94_MPORT_222_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [2047:0] hi_lo = {_WIRE_128_95,_WIRE_128_94,_WIRE_128_93,_WIRE_128_92,_WIRE_128_91,_WIRE_128_90,_WIRE_128_89,
    _WIRE_128_88,hi_lo_hi_lo,hi_lo_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_97 = tensorFile_97_MPORT_225_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_96 = tensorFile_96_MPORT_224_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_99 = tensorFile_99_MPORT_227_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_98 = tensorFile_98_MPORT_226_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_101 = tensorFile_101_MPORT_229_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_100 = tensorFile_100_MPORT_228_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_103 = tensorFile_103_MPORT_231_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_102 = tensorFile_102_MPORT_230_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [511:0] hi_hi_lo_lo = {_WIRE_128_103,_WIRE_128_102,_WIRE_128_101,_WIRE_128_100,_WIRE_128_99,_WIRE_128_98,
    _WIRE_128_97,_WIRE_128_96}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_105 = tensorFile_105_MPORT_233_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_104 = tensorFile_104_MPORT_232_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_107 = tensorFile_107_MPORT_235_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_106 = tensorFile_106_MPORT_234_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_109 = tensorFile_109_MPORT_237_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_108 = tensorFile_108_MPORT_236_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_111 = tensorFile_111_MPORT_239_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_110 = tensorFile_110_MPORT_238_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [1023:0] hi_hi_lo = {_WIRE_128_111,_WIRE_128_110,_WIRE_128_109,_WIRE_128_108,_WIRE_128_107,_WIRE_128_106,
    _WIRE_128_105,_WIRE_128_104,hi_hi_lo_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_113 = tensorFile_113_MPORT_241_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_112 = tensorFile_112_MPORT_240_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_115 = tensorFile_115_MPORT_243_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_114 = tensorFile_114_MPORT_242_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_117 = tensorFile_117_MPORT_245_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_116 = tensorFile_116_MPORT_244_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_119 = tensorFile_119_MPORT_247_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_118 = tensorFile_118_MPORT_246_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [511:0] hi_hi_hi_lo = {_WIRE_128_119,_WIRE_128_118,_WIRE_128_117,_WIRE_128_116,_WIRE_128_115,_WIRE_128_114,
    _WIRE_128_113,_WIRE_128_112}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_128_121 = tensorFile_121_MPORT_249_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_120 = tensorFile_120_MPORT_248_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_123 = tensorFile_123_MPORT_251_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_122 = tensorFile_122_MPORT_250_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_125 = tensorFile_125_MPORT_253_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_124 = tensorFile_124_MPORT_252_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_127 = tensorFile_127_MPORT_255_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [63:0] _WIRE_128_126 = tensorFile_126_MPORT_254_data; // @[TensorLoadNarrowVME.scala 284:14 TensorLoadNarrowVME.scala 284:14]
  wire [2047:0] hi_hi = {_WIRE_128_127,_WIRE_128_126,_WIRE_128_125,_WIRE_128_124,_WIRE_128_123,_WIRE_128_122,
    _WIRE_128_121,_WIRE_128_120,hi_hi_hi_lo,hi_hi_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [8191:0] _T_276 = {hi_hi,hi_lo,lo_hi,lo_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  GenVMECmd_1 vmeCmd ( // @[TensorLoadNarrowVME.scala 75:23]
    .clock(vmeCmd_clock),
    .reset(vmeCmd_reset),
    .io_start(vmeCmd_io_start),
    .io_isBusy(vmeCmd_io_isBusy),
    .io_inst(vmeCmd_io_inst),
    .io_baddr(vmeCmd_io_baddr),
    .io_vmeCmd_ready(vmeCmd_io_vmeCmd_ready),
    .io_vmeCmd_valid(vmeCmd_io_vmeCmd_valid),
    .io_vmeCmd_bits_addr(vmeCmd_io_vmeCmd_bits_addr),
    .io_vmeCmd_bits_len(vmeCmd_io_vmeCmd_bits_len),
    .io_vmeCmd_bits_tag(vmeCmd_io_vmeCmd_bits_tag),
    .io_readLen(vmeCmd_io_readLen),
    .io_done(vmeCmd_io_done)
  );
  ReadVMEData_1 readData ( // @[TensorLoadNarrowVME.scala 105:24]
    .clock(readData_clock),
    .reset(readData_reset),
    .io_start(readData_io_start),
    .io_vmeData_ready(readData_io_vmeData_ready),
    .io_vmeData_valid(readData_io_vmeData_valid),
    .io_vmeData_bits_tag(readData_io_vmeData_bits_tag),
    .io_idx(readData_io_idx),
    .io_col(readData_io_col)
  );
  ZeroPadding_1 fillPadding ( // @[TensorLoadNarrowVME.scala 119:27]
    .clock(fillPadding_clock),
    .reset(fillPadding_reset),
    .io_canWriteMem(fillPadding_io_canWriteMem),
    .io_inst(fillPadding_io_inst),
    .io_tensorIdx_valid(fillPadding_io_tensorIdx_valid),
    .io_tensorIdx_bits(fillPadding_io_tensorIdx_bits),
    .io_start(fillPadding_io_start),
    .io_done(fillPadding_io_done)
  );
  assign tensorFile_0_MPORT_128_addr = tensorFile_0_MPORT_128_addr_pipe_0;
  assign tensorFile_0_MPORT_128_data = tensorFile_0[tensorFile_0_MPORT_128_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_0_MPORT_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_0_MPORT_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_0_MPORT_mask = 1'h1;
  assign tensorFile_0_MPORT_en = _waddr_0_T ? 1'h0 : wenTensInstr_0;
  assign tensorFile_1_MPORT_129_addr = tensorFile_1_MPORT_129_addr_pipe_0;
  assign tensorFile_1_MPORT_129_data = tensorFile_1[tensorFile_1_MPORT_129_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_1_MPORT_1_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_1_MPORT_1_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_1_MPORT_1_mask = 1'h1;
  assign tensorFile_1_MPORT_1_en = _waddr_0_T ? 1'h0 : wenTensInstr_1;
  assign tensorFile_2_MPORT_130_addr = tensorFile_2_MPORT_130_addr_pipe_0;
  assign tensorFile_2_MPORT_130_data = tensorFile_2[tensorFile_2_MPORT_130_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_2_MPORT_2_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_2_MPORT_2_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_2_MPORT_2_mask = 1'h1;
  assign tensorFile_2_MPORT_2_en = _waddr_0_T ? 1'h0 : wenTensInstr_2;
  assign tensorFile_3_MPORT_131_addr = tensorFile_3_MPORT_131_addr_pipe_0;
  assign tensorFile_3_MPORT_131_data = tensorFile_3[tensorFile_3_MPORT_131_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_3_MPORT_3_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_3_MPORT_3_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_3_MPORT_3_mask = 1'h1;
  assign tensorFile_3_MPORT_3_en = _waddr_0_T ? 1'h0 : wenTensInstr_3;
  assign tensorFile_4_MPORT_132_addr = tensorFile_4_MPORT_132_addr_pipe_0;
  assign tensorFile_4_MPORT_132_data = tensorFile_4[tensorFile_4_MPORT_132_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_4_MPORT_4_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_4_MPORT_4_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_4_MPORT_4_mask = 1'h1;
  assign tensorFile_4_MPORT_4_en = _waddr_0_T ? 1'h0 : wenTensInstr_4;
  assign tensorFile_5_MPORT_133_addr = tensorFile_5_MPORT_133_addr_pipe_0;
  assign tensorFile_5_MPORT_133_data = tensorFile_5[tensorFile_5_MPORT_133_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_5_MPORT_5_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_5_MPORT_5_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_5_MPORT_5_mask = 1'h1;
  assign tensorFile_5_MPORT_5_en = _waddr_0_T ? 1'h0 : wenTensInstr_5;
  assign tensorFile_6_MPORT_134_addr = tensorFile_6_MPORT_134_addr_pipe_0;
  assign tensorFile_6_MPORT_134_data = tensorFile_6[tensorFile_6_MPORT_134_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_6_MPORT_6_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_6_MPORT_6_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_6_MPORT_6_mask = 1'h1;
  assign tensorFile_6_MPORT_6_en = _waddr_0_T ? 1'h0 : wenTensInstr_6;
  assign tensorFile_7_MPORT_135_addr = tensorFile_7_MPORT_135_addr_pipe_0;
  assign tensorFile_7_MPORT_135_data = tensorFile_7[tensorFile_7_MPORT_135_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_7_MPORT_7_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_7_MPORT_7_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_7_MPORT_7_mask = 1'h1;
  assign tensorFile_7_MPORT_7_en = _waddr_0_T ? 1'h0 : wenTensInstr_7;
  assign tensorFile_8_MPORT_136_addr = tensorFile_8_MPORT_136_addr_pipe_0;
  assign tensorFile_8_MPORT_136_data = tensorFile_8[tensorFile_8_MPORT_136_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_8_MPORT_8_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_8_MPORT_8_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_8_MPORT_8_mask = 1'h1;
  assign tensorFile_8_MPORT_8_en = _waddr_0_T ? 1'h0 : wenTensInstr_8;
  assign tensorFile_9_MPORT_137_addr = tensorFile_9_MPORT_137_addr_pipe_0;
  assign tensorFile_9_MPORT_137_data = tensorFile_9[tensorFile_9_MPORT_137_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_9_MPORT_9_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_9_MPORT_9_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_9_MPORT_9_mask = 1'h1;
  assign tensorFile_9_MPORT_9_en = _waddr_0_T ? 1'h0 : wenTensInstr_9;
  assign tensorFile_10_MPORT_138_addr = tensorFile_10_MPORT_138_addr_pipe_0;
  assign tensorFile_10_MPORT_138_data = tensorFile_10[tensorFile_10_MPORT_138_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_10_MPORT_10_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_10_MPORT_10_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_10_MPORT_10_mask = 1'h1;
  assign tensorFile_10_MPORT_10_en = _waddr_0_T ? 1'h0 : wenTensInstr_10;
  assign tensorFile_11_MPORT_139_addr = tensorFile_11_MPORT_139_addr_pipe_0;
  assign tensorFile_11_MPORT_139_data = tensorFile_11[tensorFile_11_MPORT_139_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_11_MPORT_11_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_11_MPORT_11_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_11_MPORT_11_mask = 1'h1;
  assign tensorFile_11_MPORT_11_en = _waddr_0_T ? 1'h0 : wenTensInstr_11;
  assign tensorFile_12_MPORT_140_addr = tensorFile_12_MPORT_140_addr_pipe_0;
  assign tensorFile_12_MPORT_140_data = tensorFile_12[tensorFile_12_MPORT_140_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_12_MPORT_12_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_12_MPORT_12_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_12_MPORT_12_mask = 1'h1;
  assign tensorFile_12_MPORT_12_en = _waddr_0_T ? 1'h0 : wenTensInstr_12;
  assign tensorFile_13_MPORT_141_addr = tensorFile_13_MPORT_141_addr_pipe_0;
  assign tensorFile_13_MPORT_141_data = tensorFile_13[tensorFile_13_MPORT_141_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_13_MPORT_13_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_13_MPORT_13_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_13_MPORT_13_mask = 1'h1;
  assign tensorFile_13_MPORT_13_en = _waddr_0_T ? 1'h0 : wenTensInstr_13;
  assign tensorFile_14_MPORT_142_addr = tensorFile_14_MPORT_142_addr_pipe_0;
  assign tensorFile_14_MPORT_142_data = tensorFile_14[tensorFile_14_MPORT_142_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_14_MPORT_14_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_14_MPORT_14_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_14_MPORT_14_mask = 1'h1;
  assign tensorFile_14_MPORT_14_en = _waddr_0_T ? 1'h0 : wenTensInstr_14;
  assign tensorFile_15_MPORT_143_addr = tensorFile_15_MPORT_143_addr_pipe_0;
  assign tensorFile_15_MPORT_143_data = tensorFile_15[tensorFile_15_MPORT_143_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_15_MPORT_15_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_15_MPORT_15_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_15_MPORT_15_mask = 1'h1;
  assign tensorFile_15_MPORT_15_en = _waddr_0_T ? 1'h0 : wenTensInstr_15;
  assign tensorFile_16_MPORT_144_addr = tensorFile_16_MPORT_144_addr_pipe_0;
  assign tensorFile_16_MPORT_144_data = tensorFile_16[tensorFile_16_MPORT_144_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_16_MPORT_16_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_16_MPORT_16_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_16_MPORT_16_mask = 1'h1;
  assign tensorFile_16_MPORT_16_en = _waddr_0_T ? 1'h0 : wenTensInstr_16;
  assign tensorFile_17_MPORT_145_addr = tensorFile_17_MPORT_145_addr_pipe_0;
  assign tensorFile_17_MPORT_145_data = tensorFile_17[tensorFile_17_MPORT_145_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_17_MPORT_17_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_17_MPORT_17_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_17_MPORT_17_mask = 1'h1;
  assign tensorFile_17_MPORT_17_en = _waddr_0_T ? 1'h0 : wenTensInstr_17;
  assign tensorFile_18_MPORT_146_addr = tensorFile_18_MPORT_146_addr_pipe_0;
  assign tensorFile_18_MPORT_146_data = tensorFile_18[tensorFile_18_MPORT_146_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_18_MPORT_18_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_18_MPORT_18_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_18_MPORT_18_mask = 1'h1;
  assign tensorFile_18_MPORT_18_en = _waddr_0_T ? 1'h0 : wenTensInstr_18;
  assign tensorFile_19_MPORT_147_addr = tensorFile_19_MPORT_147_addr_pipe_0;
  assign tensorFile_19_MPORT_147_data = tensorFile_19[tensorFile_19_MPORT_147_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_19_MPORT_19_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_19_MPORT_19_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_19_MPORT_19_mask = 1'h1;
  assign tensorFile_19_MPORT_19_en = _waddr_0_T ? 1'h0 : wenTensInstr_19;
  assign tensorFile_20_MPORT_148_addr = tensorFile_20_MPORT_148_addr_pipe_0;
  assign tensorFile_20_MPORT_148_data = tensorFile_20[tensorFile_20_MPORT_148_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_20_MPORT_20_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_20_MPORT_20_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_20_MPORT_20_mask = 1'h1;
  assign tensorFile_20_MPORT_20_en = _waddr_0_T ? 1'h0 : wenTensInstr_20;
  assign tensorFile_21_MPORT_149_addr = tensorFile_21_MPORT_149_addr_pipe_0;
  assign tensorFile_21_MPORT_149_data = tensorFile_21[tensorFile_21_MPORT_149_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_21_MPORT_21_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_21_MPORT_21_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_21_MPORT_21_mask = 1'h1;
  assign tensorFile_21_MPORT_21_en = _waddr_0_T ? 1'h0 : wenTensInstr_21;
  assign tensorFile_22_MPORT_150_addr = tensorFile_22_MPORT_150_addr_pipe_0;
  assign tensorFile_22_MPORT_150_data = tensorFile_22[tensorFile_22_MPORT_150_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_22_MPORT_22_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_22_MPORT_22_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_22_MPORT_22_mask = 1'h1;
  assign tensorFile_22_MPORT_22_en = _waddr_0_T ? 1'h0 : wenTensInstr_22;
  assign tensorFile_23_MPORT_151_addr = tensorFile_23_MPORT_151_addr_pipe_0;
  assign tensorFile_23_MPORT_151_data = tensorFile_23[tensorFile_23_MPORT_151_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_23_MPORT_23_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_23_MPORT_23_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_23_MPORT_23_mask = 1'h1;
  assign tensorFile_23_MPORT_23_en = _waddr_0_T ? 1'h0 : wenTensInstr_23;
  assign tensorFile_24_MPORT_152_addr = tensorFile_24_MPORT_152_addr_pipe_0;
  assign tensorFile_24_MPORT_152_data = tensorFile_24[tensorFile_24_MPORT_152_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_24_MPORT_24_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_24_MPORT_24_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_24_MPORT_24_mask = 1'h1;
  assign tensorFile_24_MPORT_24_en = _waddr_0_T ? 1'h0 : wenTensInstr_24;
  assign tensorFile_25_MPORT_153_addr = tensorFile_25_MPORT_153_addr_pipe_0;
  assign tensorFile_25_MPORT_153_data = tensorFile_25[tensorFile_25_MPORT_153_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_25_MPORT_25_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_25_MPORT_25_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_25_MPORT_25_mask = 1'h1;
  assign tensorFile_25_MPORT_25_en = _waddr_0_T ? 1'h0 : wenTensInstr_25;
  assign tensorFile_26_MPORT_154_addr = tensorFile_26_MPORT_154_addr_pipe_0;
  assign tensorFile_26_MPORT_154_data = tensorFile_26[tensorFile_26_MPORT_154_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_26_MPORT_26_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_26_MPORT_26_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_26_MPORT_26_mask = 1'h1;
  assign tensorFile_26_MPORT_26_en = _waddr_0_T ? 1'h0 : wenTensInstr_26;
  assign tensorFile_27_MPORT_155_addr = tensorFile_27_MPORT_155_addr_pipe_0;
  assign tensorFile_27_MPORT_155_data = tensorFile_27[tensorFile_27_MPORT_155_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_27_MPORT_27_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_27_MPORT_27_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_27_MPORT_27_mask = 1'h1;
  assign tensorFile_27_MPORT_27_en = _waddr_0_T ? 1'h0 : wenTensInstr_27;
  assign tensorFile_28_MPORT_156_addr = tensorFile_28_MPORT_156_addr_pipe_0;
  assign tensorFile_28_MPORT_156_data = tensorFile_28[tensorFile_28_MPORT_156_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_28_MPORT_28_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_28_MPORT_28_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_28_MPORT_28_mask = 1'h1;
  assign tensorFile_28_MPORT_28_en = _waddr_0_T ? 1'h0 : wenTensInstr_28;
  assign tensorFile_29_MPORT_157_addr = tensorFile_29_MPORT_157_addr_pipe_0;
  assign tensorFile_29_MPORT_157_data = tensorFile_29[tensorFile_29_MPORT_157_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_29_MPORT_29_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_29_MPORT_29_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_29_MPORT_29_mask = 1'h1;
  assign tensorFile_29_MPORT_29_en = _waddr_0_T ? 1'h0 : wenTensInstr_29;
  assign tensorFile_30_MPORT_158_addr = tensorFile_30_MPORT_158_addr_pipe_0;
  assign tensorFile_30_MPORT_158_data = tensorFile_30[tensorFile_30_MPORT_158_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_30_MPORT_30_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_30_MPORT_30_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_30_MPORT_30_mask = 1'h1;
  assign tensorFile_30_MPORT_30_en = _waddr_0_T ? 1'h0 : wenTensInstr_30;
  assign tensorFile_31_MPORT_159_addr = tensorFile_31_MPORT_159_addr_pipe_0;
  assign tensorFile_31_MPORT_159_data = tensorFile_31[tensorFile_31_MPORT_159_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_31_MPORT_31_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_31_MPORT_31_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_31_MPORT_31_mask = 1'h1;
  assign tensorFile_31_MPORT_31_en = _waddr_0_T ? 1'h0 : wenTensInstr_31;
  assign tensorFile_32_MPORT_160_addr = tensorFile_32_MPORT_160_addr_pipe_0;
  assign tensorFile_32_MPORT_160_data = tensorFile_32[tensorFile_32_MPORT_160_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_32_MPORT_32_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_32_MPORT_32_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_32_MPORT_32_mask = 1'h1;
  assign tensorFile_32_MPORT_32_en = _waddr_0_T ? 1'h0 : wenTensInstr_32;
  assign tensorFile_33_MPORT_161_addr = tensorFile_33_MPORT_161_addr_pipe_0;
  assign tensorFile_33_MPORT_161_data = tensorFile_33[tensorFile_33_MPORT_161_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_33_MPORT_33_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_33_MPORT_33_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_33_MPORT_33_mask = 1'h1;
  assign tensorFile_33_MPORT_33_en = _waddr_0_T ? 1'h0 : wenTensInstr_33;
  assign tensorFile_34_MPORT_162_addr = tensorFile_34_MPORT_162_addr_pipe_0;
  assign tensorFile_34_MPORT_162_data = tensorFile_34[tensorFile_34_MPORT_162_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_34_MPORT_34_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_34_MPORT_34_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_34_MPORT_34_mask = 1'h1;
  assign tensorFile_34_MPORT_34_en = _waddr_0_T ? 1'h0 : wenTensInstr_34;
  assign tensorFile_35_MPORT_163_addr = tensorFile_35_MPORT_163_addr_pipe_0;
  assign tensorFile_35_MPORT_163_data = tensorFile_35[tensorFile_35_MPORT_163_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_35_MPORT_35_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_35_MPORT_35_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_35_MPORT_35_mask = 1'h1;
  assign tensorFile_35_MPORT_35_en = _waddr_0_T ? 1'h0 : wenTensInstr_35;
  assign tensorFile_36_MPORT_164_addr = tensorFile_36_MPORT_164_addr_pipe_0;
  assign tensorFile_36_MPORT_164_data = tensorFile_36[tensorFile_36_MPORT_164_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_36_MPORT_36_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_36_MPORT_36_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_36_MPORT_36_mask = 1'h1;
  assign tensorFile_36_MPORT_36_en = _waddr_0_T ? 1'h0 : wenTensInstr_36;
  assign tensorFile_37_MPORT_165_addr = tensorFile_37_MPORT_165_addr_pipe_0;
  assign tensorFile_37_MPORT_165_data = tensorFile_37[tensorFile_37_MPORT_165_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_37_MPORT_37_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_37_MPORT_37_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_37_MPORT_37_mask = 1'h1;
  assign tensorFile_37_MPORT_37_en = _waddr_0_T ? 1'h0 : wenTensInstr_37;
  assign tensorFile_38_MPORT_166_addr = tensorFile_38_MPORT_166_addr_pipe_0;
  assign tensorFile_38_MPORT_166_data = tensorFile_38[tensorFile_38_MPORT_166_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_38_MPORT_38_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_38_MPORT_38_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_38_MPORT_38_mask = 1'h1;
  assign tensorFile_38_MPORT_38_en = _waddr_0_T ? 1'h0 : wenTensInstr_38;
  assign tensorFile_39_MPORT_167_addr = tensorFile_39_MPORT_167_addr_pipe_0;
  assign tensorFile_39_MPORT_167_data = tensorFile_39[tensorFile_39_MPORT_167_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_39_MPORT_39_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_39_MPORT_39_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_39_MPORT_39_mask = 1'h1;
  assign tensorFile_39_MPORT_39_en = _waddr_0_T ? 1'h0 : wenTensInstr_39;
  assign tensorFile_40_MPORT_168_addr = tensorFile_40_MPORT_168_addr_pipe_0;
  assign tensorFile_40_MPORT_168_data = tensorFile_40[tensorFile_40_MPORT_168_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_40_MPORT_40_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_40_MPORT_40_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_40_MPORT_40_mask = 1'h1;
  assign tensorFile_40_MPORT_40_en = _waddr_0_T ? 1'h0 : wenTensInstr_40;
  assign tensorFile_41_MPORT_169_addr = tensorFile_41_MPORT_169_addr_pipe_0;
  assign tensorFile_41_MPORT_169_data = tensorFile_41[tensorFile_41_MPORT_169_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_41_MPORT_41_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_41_MPORT_41_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_41_MPORT_41_mask = 1'h1;
  assign tensorFile_41_MPORT_41_en = _waddr_0_T ? 1'h0 : wenTensInstr_41;
  assign tensorFile_42_MPORT_170_addr = tensorFile_42_MPORT_170_addr_pipe_0;
  assign tensorFile_42_MPORT_170_data = tensorFile_42[tensorFile_42_MPORT_170_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_42_MPORT_42_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_42_MPORT_42_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_42_MPORT_42_mask = 1'h1;
  assign tensorFile_42_MPORT_42_en = _waddr_0_T ? 1'h0 : wenTensInstr_42;
  assign tensorFile_43_MPORT_171_addr = tensorFile_43_MPORT_171_addr_pipe_0;
  assign tensorFile_43_MPORT_171_data = tensorFile_43[tensorFile_43_MPORT_171_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_43_MPORT_43_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_43_MPORT_43_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_43_MPORT_43_mask = 1'h1;
  assign tensorFile_43_MPORT_43_en = _waddr_0_T ? 1'h0 : wenTensInstr_43;
  assign tensorFile_44_MPORT_172_addr = tensorFile_44_MPORT_172_addr_pipe_0;
  assign tensorFile_44_MPORT_172_data = tensorFile_44[tensorFile_44_MPORT_172_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_44_MPORT_44_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_44_MPORT_44_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_44_MPORT_44_mask = 1'h1;
  assign tensorFile_44_MPORT_44_en = _waddr_0_T ? 1'h0 : wenTensInstr_44;
  assign tensorFile_45_MPORT_173_addr = tensorFile_45_MPORT_173_addr_pipe_0;
  assign tensorFile_45_MPORT_173_data = tensorFile_45[tensorFile_45_MPORT_173_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_45_MPORT_45_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_45_MPORT_45_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_45_MPORT_45_mask = 1'h1;
  assign tensorFile_45_MPORT_45_en = _waddr_0_T ? 1'h0 : wenTensInstr_45;
  assign tensorFile_46_MPORT_174_addr = tensorFile_46_MPORT_174_addr_pipe_0;
  assign tensorFile_46_MPORT_174_data = tensorFile_46[tensorFile_46_MPORT_174_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_46_MPORT_46_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_46_MPORT_46_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_46_MPORT_46_mask = 1'h1;
  assign tensorFile_46_MPORT_46_en = _waddr_0_T ? 1'h0 : wenTensInstr_46;
  assign tensorFile_47_MPORT_175_addr = tensorFile_47_MPORT_175_addr_pipe_0;
  assign tensorFile_47_MPORT_175_data = tensorFile_47[tensorFile_47_MPORT_175_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_47_MPORT_47_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_47_MPORT_47_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_47_MPORT_47_mask = 1'h1;
  assign tensorFile_47_MPORT_47_en = _waddr_0_T ? 1'h0 : wenTensInstr_47;
  assign tensorFile_48_MPORT_176_addr = tensorFile_48_MPORT_176_addr_pipe_0;
  assign tensorFile_48_MPORT_176_data = tensorFile_48[tensorFile_48_MPORT_176_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_48_MPORT_48_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_48_MPORT_48_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_48_MPORT_48_mask = 1'h1;
  assign tensorFile_48_MPORT_48_en = _waddr_0_T ? 1'h0 : wenTensInstr_48;
  assign tensorFile_49_MPORT_177_addr = tensorFile_49_MPORT_177_addr_pipe_0;
  assign tensorFile_49_MPORT_177_data = tensorFile_49[tensorFile_49_MPORT_177_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_49_MPORT_49_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_49_MPORT_49_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_49_MPORT_49_mask = 1'h1;
  assign tensorFile_49_MPORT_49_en = _waddr_0_T ? 1'h0 : wenTensInstr_49;
  assign tensorFile_50_MPORT_178_addr = tensorFile_50_MPORT_178_addr_pipe_0;
  assign tensorFile_50_MPORT_178_data = tensorFile_50[tensorFile_50_MPORT_178_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_50_MPORT_50_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_50_MPORT_50_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_50_MPORT_50_mask = 1'h1;
  assign tensorFile_50_MPORT_50_en = _waddr_0_T ? 1'h0 : wenTensInstr_50;
  assign tensorFile_51_MPORT_179_addr = tensorFile_51_MPORT_179_addr_pipe_0;
  assign tensorFile_51_MPORT_179_data = tensorFile_51[tensorFile_51_MPORT_179_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_51_MPORT_51_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_51_MPORT_51_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_51_MPORT_51_mask = 1'h1;
  assign tensorFile_51_MPORT_51_en = _waddr_0_T ? 1'h0 : wenTensInstr_51;
  assign tensorFile_52_MPORT_180_addr = tensorFile_52_MPORT_180_addr_pipe_0;
  assign tensorFile_52_MPORT_180_data = tensorFile_52[tensorFile_52_MPORT_180_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_52_MPORT_52_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_52_MPORT_52_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_52_MPORT_52_mask = 1'h1;
  assign tensorFile_52_MPORT_52_en = _waddr_0_T ? 1'h0 : wenTensInstr_52;
  assign tensorFile_53_MPORT_181_addr = tensorFile_53_MPORT_181_addr_pipe_0;
  assign tensorFile_53_MPORT_181_data = tensorFile_53[tensorFile_53_MPORT_181_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_53_MPORT_53_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_53_MPORT_53_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_53_MPORT_53_mask = 1'h1;
  assign tensorFile_53_MPORT_53_en = _waddr_0_T ? 1'h0 : wenTensInstr_53;
  assign tensorFile_54_MPORT_182_addr = tensorFile_54_MPORT_182_addr_pipe_0;
  assign tensorFile_54_MPORT_182_data = tensorFile_54[tensorFile_54_MPORT_182_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_54_MPORT_54_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_54_MPORT_54_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_54_MPORT_54_mask = 1'h1;
  assign tensorFile_54_MPORT_54_en = _waddr_0_T ? 1'h0 : wenTensInstr_54;
  assign tensorFile_55_MPORT_183_addr = tensorFile_55_MPORT_183_addr_pipe_0;
  assign tensorFile_55_MPORT_183_data = tensorFile_55[tensorFile_55_MPORT_183_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_55_MPORT_55_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_55_MPORT_55_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_55_MPORT_55_mask = 1'h1;
  assign tensorFile_55_MPORT_55_en = _waddr_0_T ? 1'h0 : wenTensInstr_55;
  assign tensorFile_56_MPORT_184_addr = tensorFile_56_MPORT_184_addr_pipe_0;
  assign tensorFile_56_MPORT_184_data = tensorFile_56[tensorFile_56_MPORT_184_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_56_MPORT_56_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_56_MPORT_56_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_56_MPORT_56_mask = 1'h1;
  assign tensorFile_56_MPORT_56_en = _waddr_0_T ? 1'h0 : wenTensInstr_56;
  assign tensorFile_57_MPORT_185_addr = tensorFile_57_MPORT_185_addr_pipe_0;
  assign tensorFile_57_MPORT_185_data = tensorFile_57[tensorFile_57_MPORT_185_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_57_MPORT_57_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_57_MPORT_57_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_57_MPORT_57_mask = 1'h1;
  assign tensorFile_57_MPORT_57_en = _waddr_0_T ? 1'h0 : wenTensInstr_57;
  assign tensorFile_58_MPORT_186_addr = tensorFile_58_MPORT_186_addr_pipe_0;
  assign tensorFile_58_MPORT_186_data = tensorFile_58[tensorFile_58_MPORT_186_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_58_MPORT_58_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_58_MPORT_58_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_58_MPORT_58_mask = 1'h1;
  assign tensorFile_58_MPORT_58_en = _waddr_0_T ? 1'h0 : wenTensInstr_58;
  assign tensorFile_59_MPORT_187_addr = tensorFile_59_MPORT_187_addr_pipe_0;
  assign tensorFile_59_MPORT_187_data = tensorFile_59[tensorFile_59_MPORT_187_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_59_MPORT_59_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_59_MPORT_59_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_59_MPORT_59_mask = 1'h1;
  assign tensorFile_59_MPORT_59_en = _waddr_0_T ? 1'h0 : wenTensInstr_59;
  assign tensorFile_60_MPORT_188_addr = tensorFile_60_MPORT_188_addr_pipe_0;
  assign tensorFile_60_MPORT_188_data = tensorFile_60[tensorFile_60_MPORT_188_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_60_MPORT_60_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_60_MPORT_60_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_60_MPORT_60_mask = 1'h1;
  assign tensorFile_60_MPORT_60_en = _waddr_0_T ? 1'h0 : wenTensInstr_60;
  assign tensorFile_61_MPORT_189_addr = tensorFile_61_MPORT_189_addr_pipe_0;
  assign tensorFile_61_MPORT_189_data = tensorFile_61[tensorFile_61_MPORT_189_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_61_MPORT_61_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_61_MPORT_61_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_61_MPORT_61_mask = 1'h1;
  assign tensorFile_61_MPORT_61_en = _waddr_0_T ? 1'h0 : wenTensInstr_61;
  assign tensorFile_62_MPORT_190_addr = tensorFile_62_MPORT_190_addr_pipe_0;
  assign tensorFile_62_MPORT_190_data = tensorFile_62[tensorFile_62_MPORT_190_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_62_MPORT_62_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_62_MPORT_62_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_62_MPORT_62_mask = 1'h1;
  assign tensorFile_62_MPORT_62_en = _waddr_0_T ? 1'h0 : wenTensInstr_62;
  assign tensorFile_63_MPORT_191_addr = tensorFile_63_MPORT_191_addr_pipe_0;
  assign tensorFile_63_MPORT_191_data = tensorFile_63[tensorFile_63_MPORT_191_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_63_MPORT_63_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_63_MPORT_63_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_63_MPORT_63_mask = 1'h1;
  assign tensorFile_63_MPORT_63_en = _waddr_0_T ? 1'h0 : wenTensInstr_63;
  assign tensorFile_64_MPORT_192_addr = tensorFile_64_MPORT_192_addr_pipe_0;
  assign tensorFile_64_MPORT_192_data = tensorFile_64[tensorFile_64_MPORT_192_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_64_MPORT_64_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_64_MPORT_64_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_64_MPORT_64_mask = 1'h1;
  assign tensorFile_64_MPORT_64_en = _waddr_0_T ? 1'h0 : wenTensInstr_64;
  assign tensorFile_65_MPORT_193_addr = tensorFile_65_MPORT_193_addr_pipe_0;
  assign tensorFile_65_MPORT_193_data = tensorFile_65[tensorFile_65_MPORT_193_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_65_MPORT_65_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_65_MPORT_65_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_65_MPORT_65_mask = 1'h1;
  assign tensorFile_65_MPORT_65_en = _waddr_0_T ? 1'h0 : wenTensInstr_65;
  assign tensorFile_66_MPORT_194_addr = tensorFile_66_MPORT_194_addr_pipe_0;
  assign tensorFile_66_MPORT_194_data = tensorFile_66[tensorFile_66_MPORT_194_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_66_MPORT_66_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_66_MPORT_66_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_66_MPORT_66_mask = 1'h1;
  assign tensorFile_66_MPORT_66_en = _waddr_0_T ? 1'h0 : wenTensInstr_66;
  assign tensorFile_67_MPORT_195_addr = tensorFile_67_MPORT_195_addr_pipe_0;
  assign tensorFile_67_MPORT_195_data = tensorFile_67[tensorFile_67_MPORT_195_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_67_MPORT_67_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_67_MPORT_67_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_67_MPORT_67_mask = 1'h1;
  assign tensorFile_67_MPORT_67_en = _waddr_0_T ? 1'h0 : wenTensInstr_67;
  assign tensorFile_68_MPORT_196_addr = tensorFile_68_MPORT_196_addr_pipe_0;
  assign tensorFile_68_MPORT_196_data = tensorFile_68[tensorFile_68_MPORT_196_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_68_MPORT_68_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_68_MPORT_68_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_68_MPORT_68_mask = 1'h1;
  assign tensorFile_68_MPORT_68_en = _waddr_0_T ? 1'h0 : wenTensInstr_68;
  assign tensorFile_69_MPORT_197_addr = tensorFile_69_MPORT_197_addr_pipe_0;
  assign tensorFile_69_MPORT_197_data = tensorFile_69[tensorFile_69_MPORT_197_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_69_MPORT_69_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_69_MPORT_69_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_69_MPORT_69_mask = 1'h1;
  assign tensorFile_69_MPORT_69_en = _waddr_0_T ? 1'h0 : wenTensInstr_69;
  assign tensorFile_70_MPORT_198_addr = tensorFile_70_MPORT_198_addr_pipe_0;
  assign tensorFile_70_MPORT_198_data = tensorFile_70[tensorFile_70_MPORT_198_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_70_MPORT_70_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_70_MPORT_70_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_70_MPORT_70_mask = 1'h1;
  assign tensorFile_70_MPORT_70_en = _waddr_0_T ? 1'h0 : wenTensInstr_70;
  assign tensorFile_71_MPORT_199_addr = tensorFile_71_MPORT_199_addr_pipe_0;
  assign tensorFile_71_MPORT_199_data = tensorFile_71[tensorFile_71_MPORT_199_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_71_MPORT_71_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_71_MPORT_71_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_71_MPORT_71_mask = 1'h1;
  assign tensorFile_71_MPORT_71_en = _waddr_0_T ? 1'h0 : wenTensInstr_71;
  assign tensorFile_72_MPORT_200_addr = tensorFile_72_MPORT_200_addr_pipe_0;
  assign tensorFile_72_MPORT_200_data = tensorFile_72[tensorFile_72_MPORT_200_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_72_MPORT_72_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_72_MPORT_72_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_72_MPORT_72_mask = 1'h1;
  assign tensorFile_72_MPORT_72_en = _waddr_0_T ? 1'h0 : wenTensInstr_72;
  assign tensorFile_73_MPORT_201_addr = tensorFile_73_MPORT_201_addr_pipe_0;
  assign tensorFile_73_MPORT_201_data = tensorFile_73[tensorFile_73_MPORT_201_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_73_MPORT_73_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_73_MPORT_73_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_73_MPORT_73_mask = 1'h1;
  assign tensorFile_73_MPORT_73_en = _waddr_0_T ? 1'h0 : wenTensInstr_73;
  assign tensorFile_74_MPORT_202_addr = tensorFile_74_MPORT_202_addr_pipe_0;
  assign tensorFile_74_MPORT_202_data = tensorFile_74[tensorFile_74_MPORT_202_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_74_MPORT_74_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_74_MPORT_74_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_74_MPORT_74_mask = 1'h1;
  assign tensorFile_74_MPORT_74_en = _waddr_0_T ? 1'h0 : wenTensInstr_74;
  assign tensorFile_75_MPORT_203_addr = tensorFile_75_MPORT_203_addr_pipe_0;
  assign tensorFile_75_MPORT_203_data = tensorFile_75[tensorFile_75_MPORT_203_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_75_MPORT_75_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_75_MPORT_75_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_75_MPORT_75_mask = 1'h1;
  assign tensorFile_75_MPORT_75_en = _waddr_0_T ? 1'h0 : wenTensInstr_75;
  assign tensorFile_76_MPORT_204_addr = tensorFile_76_MPORT_204_addr_pipe_0;
  assign tensorFile_76_MPORT_204_data = tensorFile_76[tensorFile_76_MPORT_204_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_76_MPORT_76_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_76_MPORT_76_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_76_MPORT_76_mask = 1'h1;
  assign tensorFile_76_MPORT_76_en = _waddr_0_T ? 1'h0 : wenTensInstr_76;
  assign tensorFile_77_MPORT_205_addr = tensorFile_77_MPORT_205_addr_pipe_0;
  assign tensorFile_77_MPORT_205_data = tensorFile_77[tensorFile_77_MPORT_205_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_77_MPORT_77_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_77_MPORT_77_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_77_MPORT_77_mask = 1'h1;
  assign tensorFile_77_MPORT_77_en = _waddr_0_T ? 1'h0 : wenTensInstr_77;
  assign tensorFile_78_MPORT_206_addr = tensorFile_78_MPORT_206_addr_pipe_0;
  assign tensorFile_78_MPORT_206_data = tensorFile_78[tensorFile_78_MPORT_206_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_78_MPORT_78_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_78_MPORT_78_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_78_MPORT_78_mask = 1'h1;
  assign tensorFile_78_MPORT_78_en = _waddr_0_T ? 1'h0 : wenTensInstr_78;
  assign tensorFile_79_MPORT_207_addr = tensorFile_79_MPORT_207_addr_pipe_0;
  assign tensorFile_79_MPORT_207_data = tensorFile_79[tensorFile_79_MPORT_207_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_79_MPORT_79_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_79_MPORT_79_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_79_MPORT_79_mask = 1'h1;
  assign tensorFile_79_MPORT_79_en = _waddr_0_T ? 1'h0 : wenTensInstr_79;
  assign tensorFile_80_MPORT_208_addr = tensorFile_80_MPORT_208_addr_pipe_0;
  assign tensorFile_80_MPORT_208_data = tensorFile_80[tensorFile_80_MPORT_208_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_80_MPORT_80_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_80_MPORT_80_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_80_MPORT_80_mask = 1'h1;
  assign tensorFile_80_MPORT_80_en = _waddr_0_T ? 1'h0 : wenTensInstr_80;
  assign tensorFile_81_MPORT_209_addr = tensorFile_81_MPORT_209_addr_pipe_0;
  assign tensorFile_81_MPORT_209_data = tensorFile_81[tensorFile_81_MPORT_209_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_81_MPORT_81_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_81_MPORT_81_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_81_MPORT_81_mask = 1'h1;
  assign tensorFile_81_MPORT_81_en = _waddr_0_T ? 1'h0 : wenTensInstr_81;
  assign tensorFile_82_MPORT_210_addr = tensorFile_82_MPORT_210_addr_pipe_0;
  assign tensorFile_82_MPORT_210_data = tensorFile_82[tensorFile_82_MPORT_210_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_82_MPORT_82_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_82_MPORT_82_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_82_MPORT_82_mask = 1'h1;
  assign tensorFile_82_MPORT_82_en = _waddr_0_T ? 1'h0 : wenTensInstr_82;
  assign tensorFile_83_MPORT_211_addr = tensorFile_83_MPORT_211_addr_pipe_0;
  assign tensorFile_83_MPORT_211_data = tensorFile_83[tensorFile_83_MPORT_211_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_83_MPORT_83_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_83_MPORT_83_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_83_MPORT_83_mask = 1'h1;
  assign tensorFile_83_MPORT_83_en = _waddr_0_T ? 1'h0 : wenTensInstr_83;
  assign tensorFile_84_MPORT_212_addr = tensorFile_84_MPORT_212_addr_pipe_0;
  assign tensorFile_84_MPORT_212_data = tensorFile_84[tensorFile_84_MPORT_212_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_84_MPORT_84_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_84_MPORT_84_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_84_MPORT_84_mask = 1'h1;
  assign tensorFile_84_MPORT_84_en = _waddr_0_T ? 1'h0 : wenTensInstr_84;
  assign tensorFile_85_MPORT_213_addr = tensorFile_85_MPORT_213_addr_pipe_0;
  assign tensorFile_85_MPORT_213_data = tensorFile_85[tensorFile_85_MPORT_213_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_85_MPORT_85_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_85_MPORT_85_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_85_MPORT_85_mask = 1'h1;
  assign tensorFile_85_MPORT_85_en = _waddr_0_T ? 1'h0 : wenTensInstr_85;
  assign tensorFile_86_MPORT_214_addr = tensorFile_86_MPORT_214_addr_pipe_0;
  assign tensorFile_86_MPORT_214_data = tensorFile_86[tensorFile_86_MPORT_214_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_86_MPORT_86_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_86_MPORT_86_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_86_MPORT_86_mask = 1'h1;
  assign tensorFile_86_MPORT_86_en = _waddr_0_T ? 1'h0 : wenTensInstr_86;
  assign tensorFile_87_MPORT_215_addr = tensorFile_87_MPORT_215_addr_pipe_0;
  assign tensorFile_87_MPORT_215_data = tensorFile_87[tensorFile_87_MPORT_215_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_87_MPORT_87_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_87_MPORT_87_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_87_MPORT_87_mask = 1'h1;
  assign tensorFile_87_MPORT_87_en = _waddr_0_T ? 1'h0 : wenTensInstr_87;
  assign tensorFile_88_MPORT_216_addr = tensorFile_88_MPORT_216_addr_pipe_0;
  assign tensorFile_88_MPORT_216_data = tensorFile_88[tensorFile_88_MPORT_216_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_88_MPORT_88_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_88_MPORT_88_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_88_MPORT_88_mask = 1'h1;
  assign tensorFile_88_MPORT_88_en = _waddr_0_T ? 1'h0 : wenTensInstr_88;
  assign tensorFile_89_MPORT_217_addr = tensorFile_89_MPORT_217_addr_pipe_0;
  assign tensorFile_89_MPORT_217_data = tensorFile_89[tensorFile_89_MPORT_217_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_89_MPORT_89_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_89_MPORT_89_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_89_MPORT_89_mask = 1'h1;
  assign tensorFile_89_MPORT_89_en = _waddr_0_T ? 1'h0 : wenTensInstr_89;
  assign tensorFile_90_MPORT_218_addr = tensorFile_90_MPORT_218_addr_pipe_0;
  assign tensorFile_90_MPORT_218_data = tensorFile_90[tensorFile_90_MPORT_218_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_90_MPORT_90_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_90_MPORT_90_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_90_MPORT_90_mask = 1'h1;
  assign tensorFile_90_MPORT_90_en = _waddr_0_T ? 1'h0 : wenTensInstr_90;
  assign tensorFile_91_MPORT_219_addr = tensorFile_91_MPORT_219_addr_pipe_0;
  assign tensorFile_91_MPORT_219_data = tensorFile_91[tensorFile_91_MPORT_219_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_91_MPORT_91_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_91_MPORT_91_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_91_MPORT_91_mask = 1'h1;
  assign tensorFile_91_MPORT_91_en = _waddr_0_T ? 1'h0 : wenTensInstr_91;
  assign tensorFile_92_MPORT_220_addr = tensorFile_92_MPORT_220_addr_pipe_0;
  assign tensorFile_92_MPORT_220_data = tensorFile_92[tensorFile_92_MPORT_220_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_92_MPORT_92_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_92_MPORT_92_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_92_MPORT_92_mask = 1'h1;
  assign tensorFile_92_MPORT_92_en = _waddr_0_T ? 1'h0 : wenTensInstr_92;
  assign tensorFile_93_MPORT_221_addr = tensorFile_93_MPORT_221_addr_pipe_0;
  assign tensorFile_93_MPORT_221_data = tensorFile_93[tensorFile_93_MPORT_221_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_93_MPORT_93_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_93_MPORT_93_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_93_MPORT_93_mask = 1'h1;
  assign tensorFile_93_MPORT_93_en = _waddr_0_T ? 1'h0 : wenTensInstr_93;
  assign tensorFile_94_MPORT_222_addr = tensorFile_94_MPORT_222_addr_pipe_0;
  assign tensorFile_94_MPORT_222_data = tensorFile_94[tensorFile_94_MPORT_222_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_94_MPORT_94_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_94_MPORT_94_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_94_MPORT_94_mask = 1'h1;
  assign tensorFile_94_MPORT_94_en = _waddr_0_T ? 1'h0 : wenTensInstr_94;
  assign tensorFile_95_MPORT_223_addr = tensorFile_95_MPORT_223_addr_pipe_0;
  assign tensorFile_95_MPORT_223_data = tensorFile_95[tensorFile_95_MPORT_223_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_95_MPORT_95_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_95_MPORT_95_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_95_MPORT_95_mask = 1'h1;
  assign tensorFile_95_MPORT_95_en = _waddr_0_T ? 1'h0 : wenTensInstr_95;
  assign tensorFile_96_MPORT_224_addr = tensorFile_96_MPORT_224_addr_pipe_0;
  assign tensorFile_96_MPORT_224_data = tensorFile_96[tensorFile_96_MPORT_224_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_96_MPORT_96_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_96_MPORT_96_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_96_MPORT_96_mask = 1'h1;
  assign tensorFile_96_MPORT_96_en = _waddr_0_T ? 1'h0 : wenTensInstr_96;
  assign tensorFile_97_MPORT_225_addr = tensorFile_97_MPORT_225_addr_pipe_0;
  assign tensorFile_97_MPORT_225_data = tensorFile_97[tensorFile_97_MPORT_225_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_97_MPORT_97_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_97_MPORT_97_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_97_MPORT_97_mask = 1'h1;
  assign tensorFile_97_MPORT_97_en = _waddr_0_T ? 1'h0 : wenTensInstr_97;
  assign tensorFile_98_MPORT_226_addr = tensorFile_98_MPORT_226_addr_pipe_0;
  assign tensorFile_98_MPORT_226_data = tensorFile_98[tensorFile_98_MPORT_226_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_98_MPORT_98_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_98_MPORT_98_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_98_MPORT_98_mask = 1'h1;
  assign tensorFile_98_MPORT_98_en = _waddr_0_T ? 1'h0 : wenTensInstr_98;
  assign tensorFile_99_MPORT_227_addr = tensorFile_99_MPORT_227_addr_pipe_0;
  assign tensorFile_99_MPORT_227_data = tensorFile_99[tensorFile_99_MPORT_227_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_99_MPORT_99_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_99_MPORT_99_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_99_MPORT_99_mask = 1'h1;
  assign tensorFile_99_MPORT_99_en = _waddr_0_T ? 1'h0 : wenTensInstr_99;
  assign tensorFile_100_MPORT_228_addr = tensorFile_100_MPORT_228_addr_pipe_0;
  assign tensorFile_100_MPORT_228_data = tensorFile_100[tensorFile_100_MPORT_228_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_100_MPORT_100_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_100_MPORT_100_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_100_MPORT_100_mask = 1'h1;
  assign tensorFile_100_MPORT_100_en = _waddr_0_T ? 1'h0 : wenTensInstr_100;
  assign tensorFile_101_MPORT_229_addr = tensorFile_101_MPORT_229_addr_pipe_0;
  assign tensorFile_101_MPORT_229_data = tensorFile_101[tensorFile_101_MPORT_229_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_101_MPORT_101_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_101_MPORT_101_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_101_MPORT_101_mask = 1'h1;
  assign tensorFile_101_MPORT_101_en = _waddr_0_T ? 1'h0 : wenTensInstr_101;
  assign tensorFile_102_MPORT_230_addr = tensorFile_102_MPORT_230_addr_pipe_0;
  assign tensorFile_102_MPORT_230_data = tensorFile_102[tensorFile_102_MPORT_230_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_102_MPORT_102_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_102_MPORT_102_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_102_MPORT_102_mask = 1'h1;
  assign tensorFile_102_MPORT_102_en = _waddr_0_T ? 1'h0 : wenTensInstr_102;
  assign tensorFile_103_MPORT_231_addr = tensorFile_103_MPORT_231_addr_pipe_0;
  assign tensorFile_103_MPORT_231_data = tensorFile_103[tensorFile_103_MPORT_231_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_103_MPORT_103_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_103_MPORT_103_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_103_MPORT_103_mask = 1'h1;
  assign tensorFile_103_MPORT_103_en = _waddr_0_T ? 1'h0 : wenTensInstr_103;
  assign tensorFile_104_MPORT_232_addr = tensorFile_104_MPORT_232_addr_pipe_0;
  assign tensorFile_104_MPORT_232_data = tensorFile_104[tensorFile_104_MPORT_232_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_104_MPORT_104_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_104_MPORT_104_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_104_MPORT_104_mask = 1'h1;
  assign tensorFile_104_MPORT_104_en = _waddr_0_T ? 1'h0 : wenTensInstr_104;
  assign tensorFile_105_MPORT_233_addr = tensorFile_105_MPORT_233_addr_pipe_0;
  assign tensorFile_105_MPORT_233_data = tensorFile_105[tensorFile_105_MPORT_233_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_105_MPORT_105_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_105_MPORT_105_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_105_MPORT_105_mask = 1'h1;
  assign tensorFile_105_MPORT_105_en = _waddr_0_T ? 1'h0 : wenTensInstr_105;
  assign tensorFile_106_MPORT_234_addr = tensorFile_106_MPORT_234_addr_pipe_0;
  assign tensorFile_106_MPORT_234_data = tensorFile_106[tensorFile_106_MPORT_234_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_106_MPORT_106_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_106_MPORT_106_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_106_MPORT_106_mask = 1'h1;
  assign tensorFile_106_MPORT_106_en = _waddr_0_T ? 1'h0 : wenTensInstr_106;
  assign tensorFile_107_MPORT_235_addr = tensorFile_107_MPORT_235_addr_pipe_0;
  assign tensorFile_107_MPORT_235_data = tensorFile_107[tensorFile_107_MPORT_235_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_107_MPORT_107_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_107_MPORT_107_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_107_MPORT_107_mask = 1'h1;
  assign tensorFile_107_MPORT_107_en = _waddr_0_T ? 1'h0 : wenTensInstr_107;
  assign tensorFile_108_MPORT_236_addr = tensorFile_108_MPORT_236_addr_pipe_0;
  assign tensorFile_108_MPORT_236_data = tensorFile_108[tensorFile_108_MPORT_236_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_108_MPORT_108_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_108_MPORT_108_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_108_MPORT_108_mask = 1'h1;
  assign tensorFile_108_MPORT_108_en = _waddr_0_T ? 1'h0 : wenTensInstr_108;
  assign tensorFile_109_MPORT_237_addr = tensorFile_109_MPORT_237_addr_pipe_0;
  assign tensorFile_109_MPORT_237_data = tensorFile_109[tensorFile_109_MPORT_237_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_109_MPORT_109_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_109_MPORT_109_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_109_MPORT_109_mask = 1'h1;
  assign tensorFile_109_MPORT_109_en = _waddr_0_T ? 1'h0 : wenTensInstr_109;
  assign tensorFile_110_MPORT_238_addr = tensorFile_110_MPORT_238_addr_pipe_0;
  assign tensorFile_110_MPORT_238_data = tensorFile_110[tensorFile_110_MPORT_238_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_110_MPORT_110_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_110_MPORT_110_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_110_MPORT_110_mask = 1'h1;
  assign tensorFile_110_MPORT_110_en = _waddr_0_T ? 1'h0 : wenTensInstr_110;
  assign tensorFile_111_MPORT_239_addr = tensorFile_111_MPORT_239_addr_pipe_0;
  assign tensorFile_111_MPORT_239_data = tensorFile_111[tensorFile_111_MPORT_239_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_111_MPORT_111_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_111_MPORT_111_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_111_MPORT_111_mask = 1'h1;
  assign tensorFile_111_MPORT_111_en = _waddr_0_T ? 1'h0 : wenTensInstr_111;
  assign tensorFile_112_MPORT_240_addr = tensorFile_112_MPORT_240_addr_pipe_0;
  assign tensorFile_112_MPORT_240_data = tensorFile_112[tensorFile_112_MPORT_240_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_112_MPORT_112_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_112_MPORT_112_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_112_MPORT_112_mask = 1'h1;
  assign tensorFile_112_MPORT_112_en = _waddr_0_T ? 1'h0 : wenTensInstr_112;
  assign tensorFile_113_MPORT_241_addr = tensorFile_113_MPORT_241_addr_pipe_0;
  assign tensorFile_113_MPORT_241_data = tensorFile_113[tensorFile_113_MPORT_241_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_113_MPORT_113_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_113_MPORT_113_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_113_MPORT_113_mask = 1'h1;
  assign tensorFile_113_MPORT_113_en = _waddr_0_T ? 1'h0 : wenTensInstr_113;
  assign tensorFile_114_MPORT_242_addr = tensorFile_114_MPORT_242_addr_pipe_0;
  assign tensorFile_114_MPORT_242_data = tensorFile_114[tensorFile_114_MPORT_242_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_114_MPORT_114_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_114_MPORT_114_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_114_MPORT_114_mask = 1'h1;
  assign tensorFile_114_MPORT_114_en = _waddr_0_T ? 1'h0 : wenTensInstr_114;
  assign tensorFile_115_MPORT_243_addr = tensorFile_115_MPORT_243_addr_pipe_0;
  assign tensorFile_115_MPORT_243_data = tensorFile_115[tensorFile_115_MPORT_243_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_115_MPORT_115_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_115_MPORT_115_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_115_MPORT_115_mask = 1'h1;
  assign tensorFile_115_MPORT_115_en = _waddr_0_T ? 1'h0 : wenTensInstr_115;
  assign tensorFile_116_MPORT_244_addr = tensorFile_116_MPORT_244_addr_pipe_0;
  assign tensorFile_116_MPORT_244_data = tensorFile_116[tensorFile_116_MPORT_244_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_116_MPORT_116_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_116_MPORT_116_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_116_MPORT_116_mask = 1'h1;
  assign tensorFile_116_MPORT_116_en = _waddr_0_T ? 1'h0 : wenTensInstr_116;
  assign tensorFile_117_MPORT_245_addr = tensorFile_117_MPORT_245_addr_pipe_0;
  assign tensorFile_117_MPORT_245_data = tensorFile_117[tensorFile_117_MPORT_245_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_117_MPORT_117_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_117_MPORT_117_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_117_MPORT_117_mask = 1'h1;
  assign tensorFile_117_MPORT_117_en = _waddr_0_T ? 1'h0 : wenTensInstr_117;
  assign tensorFile_118_MPORT_246_addr = tensorFile_118_MPORT_246_addr_pipe_0;
  assign tensorFile_118_MPORT_246_data = tensorFile_118[tensorFile_118_MPORT_246_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_118_MPORT_118_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_118_MPORT_118_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_118_MPORT_118_mask = 1'h1;
  assign tensorFile_118_MPORT_118_en = _waddr_0_T ? 1'h0 : wenTensInstr_118;
  assign tensorFile_119_MPORT_247_addr = tensorFile_119_MPORT_247_addr_pipe_0;
  assign tensorFile_119_MPORT_247_data = tensorFile_119[tensorFile_119_MPORT_247_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_119_MPORT_119_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_119_MPORT_119_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_119_MPORT_119_mask = 1'h1;
  assign tensorFile_119_MPORT_119_en = _waddr_0_T ? 1'h0 : wenTensInstr_119;
  assign tensorFile_120_MPORT_248_addr = tensorFile_120_MPORT_248_addr_pipe_0;
  assign tensorFile_120_MPORT_248_data = tensorFile_120[tensorFile_120_MPORT_248_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_120_MPORT_120_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_120_MPORT_120_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_120_MPORT_120_mask = 1'h1;
  assign tensorFile_120_MPORT_120_en = _waddr_0_T ? 1'h0 : wenTensInstr_120;
  assign tensorFile_121_MPORT_249_addr = tensorFile_121_MPORT_249_addr_pipe_0;
  assign tensorFile_121_MPORT_249_data = tensorFile_121[tensorFile_121_MPORT_249_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_121_MPORT_121_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_121_MPORT_121_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_121_MPORT_121_mask = 1'h1;
  assign tensorFile_121_MPORT_121_en = _waddr_0_T ? 1'h0 : wenTensInstr_121;
  assign tensorFile_122_MPORT_250_addr = tensorFile_122_MPORT_250_addr_pipe_0;
  assign tensorFile_122_MPORT_250_data = tensorFile_122[tensorFile_122_MPORT_250_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_122_MPORT_122_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_122_MPORT_122_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_122_MPORT_122_mask = 1'h1;
  assign tensorFile_122_MPORT_122_en = _waddr_0_T ? 1'h0 : wenTensInstr_122;
  assign tensorFile_123_MPORT_251_addr = tensorFile_123_MPORT_251_addr_pipe_0;
  assign tensorFile_123_MPORT_251_data = tensorFile_123[tensorFile_123_MPORT_251_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_123_MPORT_123_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_123_MPORT_123_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_123_MPORT_123_mask = 1'h1;
  assign tensorFile_123_MPORT_123_en = _waddr_0_T ? 1'h0 : wenTensInstr_123;
  assign tensorFile_124_MPORT_252_addr = tensorFile_124_MPORT_252_addr_pipe_0;
  assign tensorFile_124_MPORT_252_data = tensorFile_124[tensorFile_124_MPORT_252_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_124_MPORT_124_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_124_MPORT_124_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_124_MPORT_124_mask = 1'h1;
  assign tensorFile_124_MPORT_124_en = _waddr_0_T ? 1'h0 : wenTensInstr_124;
  assign tensorFile_125_MPORT_253_addr = tensorFile_125_MPORT_253_addr_pipe_0;
  assign tensorFile_125_MPORT_253_data = tensorFile_125[tensorFile_125_MPORT_253_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_125_MPORT_125_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_125_MPORT_125_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_125_MPORT_125_mask = 1'h1;
  assign tensorFile_125_MPORT_125_en = _waddr_0_T ? 1'h0 : wenTensInstr_125;
  assign tensorFile_126_MPORT_254_addr = tensorFile_126_MPORT_254_addr_pipe_0;
  assign tensorFile_126_MPORT_254_data = tensorFile_126[tensorFile_126_MPORT_254_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_126_MPORT_126_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_126_MPORT_126_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_126_MPORT_126_mask = 1'h1;
  assign tensorFile_126_MPORT_126_en = _waddr_0_T ? 1'h0 : wenTensInstr_126;
  assign tensorFile_127_MPORT_255_addr = tensorFile_127_MPORT_255_addr_pipe_0;
  assign tensorFile_127_MPORT_255_data = tensorFile_127[tensorFile_127_MPORT_255_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_127_MPORT_127_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_127_MPORT_127_addr = _waddr_0_T ? 10'h0 : waddrTensInstrTmp;
  assign tensorFile_127_MPORT_127_mask = 1'h1;
  assign tensorFile_127_MPORT_127_en = _waddr_0_T ? 1'h0 : wenTensInstr_127;
  assign io_done = loadDone & fillPadding_io_done; // @[TensorLoadNarrowVME.scala 293:25]
  assign io_vme_rd_cmd_valid = vmeCmd_io_vmeCmd_valid; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_addr = vmeCmd_io_vmeCmd_bits_addr; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_len = vmeCmd_io_vmeCmd_bits_len; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_tag = vmeCmd_io_vmeCmd_bits_tag; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_data_ready = 1'h1; // @[TensorLoadNarrowVME.scala 111:24]
  assign io_tensor_rd_0_data_valid = rvalid; // @[TensorLoadNarrowVME.scala 278:36]
  assign io_tensor_rd_0_data_bits_0_0 = _T_276[31:0]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_1 = _T_276[63:32]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_2 = _T_276[95:64]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_3 = _T_276[127:96]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_4 = _T_276[159:128]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_5 = _T_276[191:160]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_6 = _T_276[223:192]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_7 = _T_276[255:224]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_8 = _T_276[287:256]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_9 = _T_276[319:288]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_10 = _T_276[351:320]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_11 = _T_276[383:352]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_12 = _T_276[415:384]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_13 = _T_276[447:416]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_14 = _T_276[479:448]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_15 = _T_276[511:480]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_0 = _T_276[543:512]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_1 = _T_276[575:544]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_2 = _T_276[607:576]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_3 = _T_276[639:608]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_4 = _T_276[671:640]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_5 = _T_276[703:672]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_6 = _T_276[735:704]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_7 = _T_276[767:736]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_8 = _T_276[799:768]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_9 = _T_276[831:800]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_10 = _T_276[863:832]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_11 = _T_276[895:864]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_12 = _T_276[927:896]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_13 = _T_276[959:928]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_14 = _T_276[991:960]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_15 = _T_276[1023:992]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_0 = _T_276[1055:1024]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_1 = _T_276[1087:1056]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_2 = _T_276[1119:1088]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_3 = _T_276[1151:1120]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_4 = _T_276[1183:1152]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_5 = _T_276[1215:1184]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_6 = _T_276[1247:1216]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_7 = _T_276[1279:1248]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_8 = _T_276[1311:1280]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_9 = _T_276[1343:1312]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_10 = _T_276[1375:1344]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_11 = _T_276[1407:1376]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_12 = _T_276[1439:1408]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_13 = _T_276[1471:1440]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_14 = _T_276[1503:1472]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_15 = _T_276[1535:1504]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_0 = _T_276[1567:1536]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_1 = _T_276[1599:1568]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_2 = _T_276[1631:1600]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_3 = _T_276[1663:1632]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_4 = _T_276[1695:1664]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_5 = _T_276[1727:1696]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_6 = _T_276[1759:1728]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_7 = _T_276[1791:1760]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_8 = _T_276[1823:1792]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_9 = _T_276[1855:1824]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_10 = _T_276[1887:1856]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_11 = _T_276[1919:1888]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_12 = _T_276[1951:1920]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_13 = _T_276[1983:1952]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_14 = _T_276[2015:1984]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_15 = _T_276[2047:2016]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_0 = _T_276[2079:2048]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_1 = _T_276[2111:2080]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_2 = _T_276[2143:2112]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_3 = _T_276[2175:2144]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_4 = _T_276[2207:2176]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_5 = _T_276[2239:2208]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_6 = _T_276[2271:2240]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_7 = _T_276[2303:2272]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_8 = _T_276[2335:2304]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_9 = _T_276[2367:2336]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_10 = _T_276[2399:2368]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_11 = _T_276[2431:2400]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_12 = _T_276[2463:2432]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_13 = _T_276[2495:2464]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_14 = _T_276[2527:2496]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_15 = _T_276[2559:2528]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_0 = _T_276[2591:2560]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_1 = _T_276[2623:2592]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_2 = _T_276[2655:2624]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_3 = _T_276[2687:2656]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_4 = _T_276[2719:2688]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_5 = _T_276[2751:2720]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_6 = _T_276[2783:2752]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_7 = _T_276[2815:2784]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_8 = _T_276[2847:2816]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_9 = _T_276[2879:2848]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_10 = _T_276[2911:2880]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_11 = _T_276[2943:2912]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_12 = _T_276[2975:2944]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_13 = _T_276[3007:2976]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_14 = _T_276[3039:3008]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_15 = _T_276[3071:3040]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_0 = _T_276[3103:3072]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_1 = _T_276[3135:3104]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_2 = _T_276[3167:3136]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_3 = _T_276[3199:3168]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_4 = _T_276[3231:3200]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_5 = _T_276[3263:3232]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_6 = _T_276[3295:3264]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_7 = _T_276[3327:3296]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_8 = _T_276[3359:3328]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_9 = _T_276[3391:3360]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_10 = _T_276[3423:3392]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_11 = _T_276[3455:3424]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_12 = _T_276[3487:3456]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_13 = _T_276[3519:3488]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_14 = _T_276[3551:3520]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_15 = _T_276[3583:3552]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_0 = _T_276[3615:3584]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_1 = _T_276[3647:3616]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_2 = _T_276[3679:3648]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_3 = _T_276[3711:3680]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_4 = _T_276[3743:3712]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_5 = _T_276[3775:3744]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_6 = _T_276[3807:3776]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_7 = _T_276[3839:3808]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_8 = _T_276[3871:3840]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_9 = _T_276[3903:3872]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_10 = _T_276[3935:3904]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_11 = _T_276[3967:3936]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_12 = _T_276[3999:3968]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_13 = _T_276[4031:4000]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_14 = _T_276[4063:4032]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_15 = _T_276[4095:4064]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_0 = _T_276[4127:4096]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_1 = _T_276[4159:4128]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_2 = _T_276[4191:4160]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_3 = _T_276[4223:4192]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_4 = _T_276[4255:4224]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_5 = _T_276[4287:4256]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_6 = _T_276[4319:4288]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_7 = _T_276[4351:4320]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_8 = _T_276[4383:4352]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_9 = _T_276[4415:4384]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_10 = _T_276[4447:4416]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_11 = _T_276[4479:4448]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_12 = _T_276[4511:4480]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_13 = _T_276[4543:4512]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_14 = _T_276[4575:4544]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_15 = _T_276[4607:4576]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_0 = _T_276[4639:4608]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_1 = _T_276[4671:4640]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_2 = _T_276[4703:4672]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_3 = _T_276[4735:4704]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_4 = _T_276[4767:4736]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_5 = _T_276[4799:4768]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_6 = _T_276[4831:4800]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_7 = _T_276[4863:4832]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_8 = _T_276[4895:4864]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_9 = _T_276[4927:4896]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_10 = _T_276[4959:4928]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_11 = _T_276[4991:4960]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_12 = _T_276[5023:4992]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_13 = _T_276[5055:5024]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_14 = _T_276[5087:5056]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_15 = _T_276[5119:5088]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_0 = _T_276[5151:5120]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_1 = _T_276[5183:5152]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_2 = _T_276[5215:5184]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_3 = _T_276[5247:5216]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_4 = _T_276[5279:5248]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_5 = _T_276[5311:5280]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_6 = _T_276[5343:5312]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_7 = _T_276[5375:5344]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_8 = _T_276[5407:5376]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_9 = _T_276[5439:5408]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_10 = _T_276[5471:5440]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_11 = _T_276[5503:5472]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_12 = _T_276[5535:5504]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_13 = _T_276[5567:5536]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_14 = _T_276[5599:5568]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_15 = _T_276[5631:5600]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_0 = _T_276[5663:5632]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_1 = _T_276[5695:5664]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_2 = _T_276[5727:5696]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_3 = _T_276[5759:5728]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_4 = _T_276[5791:5760]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_5 = _T_276[5823:5792]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_6 = _T_276[5855:5824]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_7 = _T_276[5887:5856]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_8 = _T_276[5919:5888]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_9 = _T_276[5951:5920]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_10 = _T_276[5983:5952]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_11 = _T_276[6015:5984]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_12 = _T_276[6047:6016]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_13 = _T_276[6079:6048]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_14 = _T_276[6111:6080]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_15 = _T_276[6143:6112]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_0 = _T_276[6175:6144]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_1 = _T_276[6207:6176]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_2 = _T_276[6239:6208]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_3 = _T_276[6271:6240]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_4 = _T_276[6303:6272]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_5 = _T_276[6335:6304]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_6 = _T_276[6367:6336]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_7 = _T_276[6399:6368]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_8 = _T_276[6431:6400]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_9 = _T_276[6463:6432]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_10 = _T_276[6495:6464]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_11 = _T_276[6527:6496]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_12 = _T_276[6559:6528]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_13 = _T_276[6591:6560]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_14 = _T_276[6623:6592]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_15 = _T_276[6655:6624]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_0 = _T_276[6687:6656]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_1 = _T_276[6719:6688]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_2 = _T_276[6751:6720]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_3 = _T_276[6783:6752]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_4 = _T_276[6815:6784]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_5 = _T_276[6847:6816]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_6 = _T_276[6879:6848]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_7 = _T_276[6911:6880]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_8 = _T_276[6943:6912]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_9 = _T_276[6975:6944]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_10 = _T_276[7007:6976]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_11 = _T_276[7039:7008]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_12 = _T_276[7071:7040]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_13 = _T_276[7103:7072]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_14 = _T_276[7135:7104]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_15 = _T_276[7167:7136]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_0 = _T_276[7199:7168]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_1 = _T_276[7231:7200]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_2 = _T_276[7263:7232]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_3 = _T_276[7295:7264]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_4 = _T_276[7327:7296]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_5 = _T_276[7359:7328]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_6 = _T_276[7391:7360]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_7 = _T_276[7423:7392]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_8 = _T_276[7455:7424]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_9 = _T_276[7487:7456]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_10 = _T_276[7519:7488]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_11 = _T_276[7551:7520]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_12 = _T_276[7583:7552]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_13 = _T_276[7615:7584]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_14 = _T_276[7647:7616]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_15 = _T_276[7679:7648]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_0 = _T_276[7711:7680]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_1 = _T_276[7743:7712]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_2 = _T_276[7775:7744]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_3 = _T_276[7807:7776]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_4 = _T_276[7839:7808]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_5 = _T_276[7871:7840]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_6 = _T_276[7903:7872]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_7 = _T_276[7935:7904]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_8 = _T_276[7967:7936]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_9 = _T_276[7999:7968]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_10 = _T_276[8031:8000]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_11 = _T_276[8063:8032]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_12 = _T_276[8095:8064]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_13 = _T_276[8127:8096]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_14 = _T_276[8159:8128]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_15 = _T_276[8191:8160]; // @[TensorLoadNarrowVME.scala 288:18]
  assign vmeCmd_clock = clock;
  assign vmeCmd_reset = reset;
  assign vmeCmd_io_start = io_start; // @[TensorLoadNarrowVME.scala 76:19]
  assign vmeCmd_io_isBusy = state; // @[TensorLoadNarrowVME.scala 56:22]
  assign vmeCmd_io_inst = io_inst; // @[TensorLoadNarrowVME.scala 78:18]
  assign vmeCmd_io_baddr = io_baddr; // @[TensorLoadNarrowVME.scala 79:19]
  assign vmeCmd_io_vmeCmd_ready = io_vme_rd_cmd_ready; // @[TensorLoadNarrowVME.scala 80:20]
  assign readData_clock = clock;
  assign readData_reset = reset;
  assign readData_io_start = io_start; // @[TensorLoadNarrowVME.scala 106:21]
  assign readData_io_vmeData_valid = vmeDataValidPipe; // @[TensorLoadNarrowVME.scala 107:29]
  assign readData_io_vmeData_bits_tag = vmeDataBitsPipe_tag; // @[TensorLoadNarrowVME.scala 108:28]
  assign fillPadding_clock = clock;
  assign fillPadding_reset = reset;
  assign fillPadding_io_canWriteMem = ~vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 120:33]
  assign fillPadding_io_inst = fillPadding_io_inst_REG; // @[TensorLoadNarrowVME.scala 121:23]
  assign fillPadding_io_start = fillPadding_io_start_REG; // @[TensorLoadNarrowVME.scala 122:24]
  always @(posedge clock) begin
    if(tensorFile_0_MPORT_en & tensorFile_0_MPORT_mask) begin
      tensorFile_0[tensorFile_0_MPORT_addr] <= tensorFile_0_MPORT_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_0_MPORT_128_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_0_MPORT_128_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_1_MPORT_1_en & tensorFile_1_MPORT_1_mask) begin
      tensorFile_1[tensorFile_1_MPORT_1_addr] <= tensorFile_1_MPORT_1_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_1_MPORT_129_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_1_MPORT_129_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_2_MPORT_2_en & tensorFile_2_MPORT_2_mask) begin
      tensorFile_2[tensorFile_2_MPORT_2_addr] <= tensorFile_2_MPORT_2_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_2_MPORT_130_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_2_MPORT_130_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_3_MPORT_3_en & tensorFile_3_MPORT_3_mask) begin
      tensorFile_3[tensorFile_3_MPORT_3_addr] <= tensorFile_3_MPORT_3_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_3_MPORT_131_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_3_MPORT_131_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_4_MPORT_4_en & tensorFile_4_MPORT_4_mask) begin
      tensorFile_4[tensorFile_4_MPORT_4_addr] <= tensorFile_4_MPORT_4_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_4_MPORT_132_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_4_MPORT_132_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_5_MPORT_5_en & tensorFile_5_MPORT_5_mask) begin
      tensorFile_5[tensorFile_5_MPORT_5_addr] <= tensorFile_5_MPORT_5_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_5_MPORT_133_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_5_MPORT_133_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_6_MPORT_6_en & tensorFile_6_MPORT_6_mask) begin
      tensorFile_6[tensorFile_6_MPORT_6_addr] <= tensorFile_6_MPORT_6_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_6_MPORT_134_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_6_MPORT_134_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_7_MPORT_7_en & tensorFile_7_MPORT_7_mask) begin
      tensorFile_7[tensorFile_7_MPORT_7_addr] <= tensorFile_7_MPORT_7_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_7_MPORT_135_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_7_MPORT_135_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_8_MPORT_8_en & tensorFile_8_MPORT_8_mask) begin
      tensorFile_8[tensorFile_8_MPORT_8_addr] <= tensorFile_8_MPORT_8_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_8_MPORT_136_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_8_MPORT_136_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_9_MPORT_9_en & tensorFile_9_MPORT_9_mask) begin
      tensorFile_9[tensorFile_9_MPORT_9_addr] <= tensorFile_9_MPORT_9_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_9_MPORT_137_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_9_MPORT_137_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_10_MPORT_10_en & tensorFile_10_MPORT_10_mask) begin
      tensorFile_10[tensorFile_10_MPORT_10_addr] <= tensorFile_10_MPORT_10_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_10_MPORT_138_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_10_MPORT_138_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_11_MPORT_11_en & tensorFile_11_MPORT_11_mask) begin
      tensorFile_11[tensorFile_11_MPORT_11_addr] <= tensorFile_11_MPORT_11_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_11_MPORT_139_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_11_MPORT_139_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_12_MPORT_12_en & tensorFile_12_MPORT_12_mask) begin
      tensorFile_12[tensorFile_12_MPORT_12_addr] <= tensorFile_12_MPORT_12_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_12_MPORT_140_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_12_MPORT_140_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_13_MPORT_13_en & tensorFile_13_MPORT_13_mask) begin
      tensorFile_13[tensorFile_13_MPORT_13_addr] <= tensorFile_13_MPORT_13_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_13_MPORT_141_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_13_MPORT_141_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_14_MPORT_14_en & tensorFile_14_MPORT_14_mask) begin
      tensorFile_14[tensorFile_14_MPORT_14_addr] <= tensorFile_14_MPORT_14_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_14_MPORT_142_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_14_MPORT_142_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_15_MPORT_15_en & tensorFile_15_MPORT_15_mask) begin
      tensorFile_15[tensorFile_15_MPORT_15_addr] <= tensorFile_15_MPORT_15_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_15_MPORT_143_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_15_MPORT_143_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_16_MPORT_16_en & tensorFile_16_MPORT_16_mask) begin
      tensorFile_16[tensorFile_16_MPORT_16_addr] <= tensorFile_16_MPORT_16_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_16_MPORT_144_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_16_MPORT_144_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_17_MPORT_17_en & tensorFile_17_MPORT_17_mask) begin
      tensorFile_17[tensorFile_17_MPORT_17_addr] <= tensorFile_17_MPORT_17_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_17_MPORT_145_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_17_MPORT_145_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_18_MPORT_18_en & tensorFile_18_MPORT_18_mask) begin
      tensorFile_18[tensorFile_18_MPORT_18_addr] <= tensorFile_18_MPORT_18_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_18_MPORT_146_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_18_MPORT_146_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_19_MPORT_19_en & tensorFile_19_MPORT_19_mask) begin
      tensorFile_19[tensorFile_19_MPORT_19_addr] <= tensorFile_19_MPORT_19_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_19_MPORT_147_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_19_MPORT_147_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_20_MPORT_20_en & tensorFile_20_MPORT_20_mask) begin
      tensorFile_20[tensorFile_20_MPORT_20_addr] <= tensorFile_20_MPORT_20_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_20_MPORT_148_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_20_MPORT_148_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_21_MPORT_21_en & tensorFile_21_MPORT_21_mask) begin
      tensorFile_21[tensorFile_21_MPORT_21_addr] <= tensorFile_21_MPORT_21_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_21_MPORT_149_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_21_MPORT_149_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_22_MPORT_22_en & tensorFile_22_MPORT_22_mask) begin
      tensorFile_22[tensorFile_22_MPORT_22_addr] <= tensorFile_22_MPORT_22_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_22_MPORT_150_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_22_MPORT_150_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_23_MPORT_23_en & tensorFile_23_MPORT_23_mask) begin
      tensorFile_23[tensorFile_23_MPORT_23_addr] <= tensorFile_23_MPORT_23_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_23_MPORT_151_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_23_MPORT_151_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_24_MPORT_24_en & tensorFile_24_MPORT_24_mask) begin
      tensorFile_24[tensorFile_24_MPORT_24_addr] <= tensorFile_24_MPORT_24_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_24_MPORT_152_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_24_MPORT_152_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_25_MPORT_25_en & tensorFile_25_MPORT_25_mask) begin
      tensorFile_25[tensorFile_25_MPORT_25_addr] <= tensorFile_25_MPORT_25_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_25_MPORT_153_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_25_MPORT_153_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_26_MPORT_26_en & tensorFile_26_MPORT_26_mask) begin
      tensorFile_26[tensorFile_26_MPORT_26_addr] <= tensorFile_26_MPORT_26_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_26_MPORT_154_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_26_MPORT_154_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_27_MPORT_27_en & tensorFile_27_MPORT_27_mask) begin
      tensorFile_27[tensorFile_27_MPORT_27_addr] <= tensorFile_27_MPORT_27_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_27_MPORT_155_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_27_MPORT_155_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_28_MPORT_28_en & tensorFile_28_MPORT_28_mask) begin
      tensorFile_28[tensorFile_28_MPORT_28_addr] <= tensorFile_28_MPORT_28_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_28_MPORT_156_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_28_MPORT_156_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_29_MPORT_29_en & tensorFile_29_MPORT_29_mask) begin
      tensorFile_29[tensorFile_29_MPORT_29_addr] <= tensorFile_29_MPORT_29_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_29_MPORT_157_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_29_MPORT_157_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_30_MPORT_30_en & tensorFile_30_MPORT_30_mask) begin
      tensorFile_30[tensorFile_30_MPORT_30_addr] <= tensorFile_30_MPORT_30_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_30_MPORT_158_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_30_MPORT_158_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_31_MPORT_31_en & tensorFile_31_MPORT_31_mask) begin
      tensorFile_31[tensorFile_31_MPORT_31_addr] <= tensorFile_31_MPORT_31_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_31_MPORT_159_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_31_MPORT_159_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_32_MPORT_32_en & tensorFile_32_MPORT_32_mask) begin
      tensorFile_32[tensorFile_32_MPORT_32_addr] <= tensorFile_32_MPORT_32_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_32_MPORT_160_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_32_MPORT_160_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_33_MPORT_33_en & tensorFile_33_MPORT_33_mask) begin
      tensorFile_33[tensorFile_33_MPORT_33_addr] <= tensorFile_33_MPORT_33_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_33_MPORT_161_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_33_MPORT_161_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_34_MPORT_34_en & tensorFile_34_MPORT_34_mask) begin
      tensorFile_34[tensorFile_34_MPORT_34_addr] <= tensorFile_34_MPORT_34_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_34_MPORT_162_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_34_MPORT_162_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_35_MPORT_35_en & tensorFile_35_MPORT_35_mask) begin
      tensorFile_35[tensorFile_35_MPORT_35_addr] <= tensorFile_35_MPORT_35_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_35_MPORT_163_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_35_MPORT_163_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_36_MPORT_36_en & tensorFile_36_MPORT_36_mask) begin
      tensorFile_36[tensorFile_36_MPORT_36_addr] <= tensorFile_36_MPORT_36_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_36_MPORT_164_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_36_MPORT_164_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_37_MPORT_37_en & tensorFile_37_MPORT_37_mask) begin
      tensorFile_37[tensorFile_37_MPORT_37_addr] <= tensorFile_37_MPORT_37_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_37_MPORT_165_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_37_MPORT_165_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_38_MPORT_38_en & tensorFile_38_MPORT_38_mask) begin
      tensorFile_38[tensorFile_38_MPORT_38_addr] <= tensorFile_38_MPORT_38_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_38_MPORT_166_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_38_MPORT_166_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_39_MPORT_39_en & tensorFile_39_MPORT_39_mask) begin
      tensorFile_39[tensorFile_39_MPORT_39_addr] <= tensorFile_39_MPORT_39_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_39_MPORT_167_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_39_MPORT_167_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_40_MPORT_40_en & tensorFile_40_MPORT_40_mask) begin
      tensorFile_40[tensorFile_40_MPORT_40_addr] <= tensorFile_40_MPORT_40_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_40_MPORT_168_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_40_MPORT_168_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_41_MPORT_41_en & tensorFile_41_MPORT_41_mask) begin
      tensorFile_41[tensorFile_41_MPORT_41_addr] <= tensorFile_41_MPORT_41_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_41_MPORT_169_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_41_MPORT_169_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_42_MPORT_42_en & tensorFile_42_MPORT_42_mask) begin
      tensorFile_42[tensorFile_42_MPORT_42_addr] <= tensorFile_42_MPORT_42_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_42_MPORT_170_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_42_MPORT_170_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_43_MPORT_43_en & tensorFile_43_MPORT_43_mask) begin
      tensorFile_43[tensorFile_43_MPORT_43_addr] <= tensorFile_43_MPORT_43_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_43_MPORT_171_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_43_MPORT_171_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_44_MPORT_44_en & tensorFile_44_MPORT_44_mask) begin
      tensorFile_44[tensorFile_44_MPORT_44_addr] <= tensorFile_44_MPORT_44_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_44_MPORT_172_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_44_MPORT_172_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_45_MPORT_45_en & tensorFile_45_MPORT_45_mask) begin
      tensorFile_45[tensorFile_45_MPORT_45_addr] <= tensorFile_45_MPORT_45_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_45_MPORT_173_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_45_MPORT_173_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_46_MPORT_46_en & tensorFile_46_MPORT_46_mask) begin
      tensorFile_46[tensorFile_46_MPORT_46_addr] <= tensorFile_46_MPORT_46_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_46_MPORT_174_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_46_MPORT_174_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_47_MPORT_47_en & tensorFile_47_MPORT_47_mask) begin
      tensorFile_47[tensorFile_47_MPORT_47_addr] <= tensorFile_47_MPORT_47_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_47_MPORT_175_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_47_MPORT_175_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_48_MPORT_48_en & tensorFile_48_MPORT_48_mask) begin
      tensorFile_48[tensorFile_48_MPORT_48_addr] <= tensorFile_48_MPORT_48_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_48_MPORT_176_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_48_MPORT_176_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_49_MPORT_49_en & tensorFile_49_MPORT_49_mask) begin
      tensorFile_49[tensorFile_49_MPORT_49_addr] <= tensorFile_49_MPORT_49_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_49_MPORT_177_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_49_MPORT_177_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_50_MPORT_50_en & tensorFile_50_MPORT_50_mask) begin
      tensorFile_50[tensorFile_50_MPORT_50_addr] <= tensorFile_50_MPORT_50_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_50_MPORT_178_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_50_MPORT_178_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_51_MPORT_51_en & tensorFile_51_MPORT_51_mask) begin
      tensorFile_51[tensorFile_51_MPORT_51_addr] <= tensorFile_51_MPORT_51_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_51_MPORT_179_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_51_MPORT_179_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_52_MPORT_52_en & tensorFile_52_MPORT_52_mask) begin
      tensorFile_52[tensorFile_52_MPORT_52_addr] <= tensorFile_52_MPORT_52_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_52_MPORT_180_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_52_MPORT_180_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_53_MPORT_53_en & tensorFile_53_MPORT_53_mask) begin
      tensorFile_53[tensorFile_53_MPORT_53_addr] <= tensorFile_53_MPORT_53_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_53_MPORT_181_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_53_MPORT_181_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_54_MPORT_54_en & tensorFile_54_MPORT_54_mask) begin
      tensorFile_54[tensorFile_54_MPORT_54_addr] <= tensorFile_54_MPORT_54_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_54_MPORT_182_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_54_MPORT_182_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_55_MPORT_55_en & tensorFile_55_MPORT_55_mask) begin
      tensorFile_55[tensorFile_55_MPORT_55_addr] <= tensorFile_55_MPORT_55_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_55_MPORT_183_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_55_MPORT_183_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_56_MPORT_56_en & tensorFile_56_MPORT_56_mask) begin
      tensorFile_56[tensorFile_56_MPORT_56_addr] <= tensorFile_56_MPORT_56_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_56_MPORT_184_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_56_MPORT_184_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_57_MPORT_57_en & tensorFile_57_MPORT_57_mask) begin
      tensorFile_57[tensorFile_57_MPORT_57_addr] <= tensorFile_57_MPORT_57_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_57_MPORT_185_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_57_MPORT_185_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_58_MPORT_58_en & tensorFile_58_MPORT_58_mask) begin
      tensorFile_58[tensorFile_58_MPORT_58_addr] <= tensorFile_58_MPORT_58_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_58_MPORT_186_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_58_MPORT_186_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_59_MPORT_59_en & tensorFile_59_MPORT_59_mask) begin
      tensorFile_59[tensorFile_59_MPORT_59_addr] <= tensorFile_59_MPORT_59_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_59_MPORT_187_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_59_MPORT_187_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_60_MPORT_60_en & tensorFile_60_MPORT_60_mask) begin
      tensorFile_60[tensorFile_60_MPORT_60_addr] <= tensorFile_60_MPORT_60_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_60_MPORT_188_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_60_MPORT_188_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_61_MPORT_61_en & tensorFile_61_MPORT_61_mask) begin
      tensorFile_61[tensorFile_61_MPORT_61_addr] <= tensorFile_61_MPORT_61_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_61_MPORT_189_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_61_MPORT_189_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_62_MPORT_62_en & tensorFile_62_MPORT_62_mask) begin
      tensorFile_62[tensorFile_62_MPORT_62_addr] <= tensorFile_62_MPORT_62_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_62_MPORT_190_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_62_MPORT_190_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_63_MPORT_63_en & tensorFile_63_MPORT_63_mask) begin
      tensorFile_63[tensorFile_63_MPORT_63_addr] <= tensorFile_63_MPORT_63_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_63_MPORT_191_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_63_MPORT_191_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_64_MPORT_64_en & tensorFile_64_MPORT_64_mask) begin
      tensorFile_64[tensorFile_64_MPORT_64_addr] <= tensorFile_64_MPORT_64_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_64_MPORT_192_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_64_MPORT_192_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_65_MPORT_65_en & tensorFile_65_MPORT_65_mask) begin
      tensorFile_65[tensorFile_65_MPORT_65_addr] <= tensorFile_65_MPORT_65_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_65_MPORT_193_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_65_MPORT_193_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_66_MPORT_66_en & tensorFile_66_MPORT_66_mask) begin
      tensorFile_66[tensorFile_66_MPORT_66_addr] <= tensorFile_66_MPORT_66_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_66_MPORT_194_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_66_MPORT_194_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_67_MPORT_67_en & tensorFile_67_MPORT_67_mask) begin
      tensorFile_67[tensorFile_67_MPORT_67_addr] <= tensorFile_67_MPORT_67_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_67_MPORT_195_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_67_MPORT_195_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_68_MPORT_68_en & tensorFile_68_MPORT_68_mask) begin
      tensorFile_68[tensorFile_68_MPORT_68_addr] <= tensorFile_68_MPORT_68_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_68_MPORT_196_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_68_MPORT_196_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_69_MPORT_69_en & tensorFile_69_MPORT_69_mask) begin
      tensorFile_69[tensorFile_69_MPORT_69_addr] <= tensorFile_69_MPORT_69_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_69_MPORT_197_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_69_MPORT_197_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_70_MPORT_70_en & tensorFile_70_MPORT_70_mask) begin
      tensorFile_70[tensorFile_70_MPORT_70_addr] <= tensorFile_70_MPORT_70_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_70_MPORT_198_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_70_MPORT_198_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_71_MPORT_71_en & tensorFile_71_MPORT_71_mask) begin
      tensorFile_71[tensorFile_71_MPORT_71_addr] <= tensorFile_71_MPORT_71_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_71_MPORT_199_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_71_MPORT_199_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_72_MPORT_72_en & tensorFile_72_MPORT_72_mask) begin
      tensorFile_72[tensorFile_72_MPORT_72_addr] <= tensorFile_72_MPORT_72_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_72_MPORT_200_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_72_MPORT_200_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_73_MPORT_73_en & tensorFile_73_MPORT_73_mask) begin
      tensorFile_73[tensorFile_73_MPORT_73_addr] <= tensorFile_73_MPORT_73_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_73_MPORT_201_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_73_MPORT_201_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_74_MPORT_74_en & tensorFile_74_MPORT_74_mask) begin
      tensorFile_74[tensorFile_74_MPORT_74_addr] <= tensorFile_74_MPORT_74_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_74_MPORT_202_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_74_MPORT_202_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_75_MPORT_75_en & tensorFile_75_MPORT_75_mask) begin
      tensorFile_75[tensorFile_75_MPORT_75_addr] <= tensorFile_75_MPORT_75_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_75_MPORT_203_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_75_MPORT_203_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_76_MPORT_76_en & tensorFile_76_MPORT_76_mask) begin
      tensorFile_76[tensorFile_76_MPORT_76_addr] <= tensorFile_76_MPORT_76_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_76_MPORT_204_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_76_MPORT_204_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_77_MPORT_77_en & tensorFile_77_MPORT_77_mask) begin
      tensorFile_77[tensorFile_77_MPORT_77_addr] <= tensorFile_77_MPORT_77_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_77_MPORT_205_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_77_MPORT_205_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_78_MPORT_78_en & tensorFile_78_MPORT_78_mask) begin
      tensorFile_78[tensorFile_78_MPORT_78_addr] <= tensorFile_78_MPORT_78_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_78_MPORT_206_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_78_MPORT_206_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_79_MPORT_79_en & tensorFile_79_MPORT_79_mask) begin
      tensorFile_79[tensorFile_79_MPORT_79_addr] <= tensorFile_79_MPORT_79_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_79_MPORT_207_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_79_MPORT_207_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_80_MPORT_80_en & tensorFile_80_MPORT_80_mask) begin
      tensorFile_80[tensorFile_80_MPORT_80_addr] <= tensorFile_80_MPORT_80_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_80_MPORT_208_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_80_MPORT_208_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_81_MPORT_81_en & tensorFile_81_MPORT_81_mask) begin
      tensorFile_81[tensorFile_81_MPORT_81_addr] <= tensorFile_81_MPORT_81_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_81_MPORT_209_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_81_MPORT_209_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_82_MPORT_82_en & tensorFile_82_MPORT_82_mask) begin
      tensorFile_82[tensorFile_82_MPORT_82_addr] <= tensorFile_82_MPORT_82_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_82_MPORT_210_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_82_MPORT_210_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_83_MPORT_83_en & tensorFile_83_MPORT_83_mask) begin
      tensorFile_83[tensorFile_83_MPORT_83_addr] <= tensorFile_83_MPORT_83_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_83_MPORT_211_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_83_MPORT_211_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_84_MPORT_84_en & tensorFile_84_MPORT_84_mask) begin
      tensorFile_84[tensorFile_84_MPORT_84_addr] <= tensorFile_84_MPORT_84_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_84_MPORT_212_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_84_MPORT_212_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_85_MPORT_85_en & tensorFile_85_MPORT_85_mask) begin
      tensorFile_85[tensorFile_85_MPORT_85_addr] <= tensorFile_85_MPORT_85_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_85_MPORT_213_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_85_MPORT_213_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_86_MPORT_86_en & tensorFile_86_MPORT_86_mask) begin
      tensorFile_86[tensorFile_86_MPORT_86_addr] <= tensorFile_86_MPORT_86_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_86_MPORT_214_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_86_MPORT_214_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_87_MPORT_87_en & tensorFile_87_MPORT_87_mask) begin
      tensorFile_87[tensorFile_87_MPORT_87_addr] <= tensorFile_87_MPORT_87_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_87_MPORT_215_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_87_MPORT_215_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_88_MPORT_88_en & tensorFile_88_MPORT_88_mask) begin
      tensorFile_88[tensorFile_88_MPORT_88_addr] <= tensorFile_88_MPORT_88_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_88_MPORT_216_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_88_MPORT_216_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_89_MPORT_89_en & tensorFile_89_MPORT_89_mask) begin
      tensorFile_89[tensorFile_89_MPORT_89_addr] <= tensorFile_89_MPORT_89_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_89_MPORT_217_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_89_MPORT_217_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_90_MPORT_90_en & tensorFile_90_MPORT_90_mask) begin
      tensorFile_90[tensorFile_90_MPORT_90_addr] <= tensorFile_90_MPORT_90_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_90_MPORT_218_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_90_MPORT_218_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_91_MPORT_91_en & tensorFile_91_MPORT_91_mask) begin
      tensorFile_91[tensorFile_91_MPORT_91_addr] <= tensorFile_91_MPORT_91_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_91_MPORT_219_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_91_MPORT_219_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_92_MPORT_92_en & tensorFile_92_MPORT_92_mask) begin
      tensorFile_92[tensorFile_92_MPORT_92_addr] <= tensorFile_92_MPORT_92_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_92_MPORT_220_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_92_MPORT_220_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_93_MPORT_93_en & tensorFile_93_MPORT_93_mask) begin
      tensorFile_93[tensorFile_93_MPORT_93_addr] <= tensorFile_93_MPORT_93_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_93_MPORT_221_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_93_MPORT_221_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_94_MPORT_94_en & tensorFile_94_MPORT_94_mask) begin
      tensorFile_94[tensorFile_94_MPORT_94_addr] <= tensorFile_94_MPORT_94_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_94_MPORT_222_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_94_MPORT_222_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_95_MPORT_95_en & tensorFile_95_MPORT_95_mask) begin
      tensorFile_95[tensorFile_95_MPORT_95_addr] <= tensorFile_95_MPORT_95_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_95_MPORT_223_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_95_MPORT_223_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_96_MPORT_96_en & tensorFile_96_MPORT_96_mask) begin
      tensorFile_96[tensorFile_96_MPORT_96_addr] <= tensorFile_96_MPORT_96_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_96_MPORT_224_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_96_MPORT_224_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_97_MPORT_97_en & tensorFile_97_MPORT_97_mask) begin
      tensorFile_97[tensorFile_97_MPORT_97_addr] <= tensorFile_97_MPORT_97_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_97_MPORT_225_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_97_MPORT_225_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_98_MPORT_98_en & tensorFile_98_MPORT_98_mask) begin
      tensorFile_98[tensorFile_98_MPORT_98_addr] <= tensorFile_98_MPORT_98_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_98_MPORT_226_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_98_MPORT_226_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_99_MPORT_99_en & tensorFile_99_MPORT_99_mask) begin
      tensorFile_99[tensorFile_99_MPORT_99_addr] <= tensorFile_99_MPORT_99_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_99_MPORT_227_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_99_MPORT_227_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_100_MPORT_100_en & tensorFile_100_MPORT_100_mask) begin
      tensorFile_100[tensorFile_100_MPORT_100_addr] <= tensorFile_100_MPORT_100_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_100_MPORT_228_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_100_MPORT_228_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_101_MPORT_101_en & tensorFile_101_MPORT_101_mask) begin
      tensorFile_101[tensorFile_101_MPORT_101_addr] <= tensorFile_101_MPORT_101_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_101_MPORT_229_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_101_MPORT_229_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_102_MPORT_102_en & tensorFile_102_MPORT_102_mask) begin
      tensorFile_102[tensorFile_102_MPORT_102_addr] <= tensorFile_102_MPORT_102_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_102_MPORT_230_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_102_MPORT_230_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_103_MPORT_103_en & tensorFile_103_MPORT_103_mask) begin
      tensorFile_103[tensorFile_103_MPORT_103_addr] <= tensorFile_103_MPORT_103_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_103_MPORT_231_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_103_MPORT_231_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_104_MPORT_104_en & tensorFile_104_MPORT_104_mask) begin
      tensorFile_104[tensorFile_104_MPORT_104_addr] <= tensorFile_104_MPORT_104_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_104_MPORT_232_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_104_MPORT_232_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_105_MPORT_105_en & tensorFile_105_MPORT_105_mask) begin
      tensorFile_105[tensorFile_105_MPORT_105_addr] <= tensorFile_105_MPORT_105_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_105_MPORT_233_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_105_MPORT_233_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_106_MPORT_106_en & tensorFile_106_MPORT_106_mask) begin
      tensorFile_106[tensorFile_106_MPORT_106_addr] <= tensorFile_106_MPORT_106_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_106_MPORT_234_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_106_MPORT_234_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_107_MPORT_107_en & tensorFile_107_MPORT_107_mask) begin
      tensorFile_107[tensorFile_107_MPORT_107_addr] <= tensorFile_107_MPORT_107_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_107_MPORT_235_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_107_MPORT_235_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_108_MPORT_108_en & tensorFile_108_MPORT_108_mask) begin
      tensorFile_108[tensorFile_108_MPORT_108_addr] <= tensorFile_108_MPORT_108_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_108_MPORT_236_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_108_MPORT_236_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_109_MPORT_109_en & tensorFile_109_MPORT_109_mask) begin
      tensorFile_109[tensorFile_109_MPORT_109_addr] <= tensorFile_109_MPORT_109_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_109_MPORT_237_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_109_MPORT_237_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_110_MPORT_110_en & tensorFile_110_MPORT_110_mask) begin
      tensorFile_110[tensorFile_110_MPORT_110_addr] <= tensorFile_110_MPORT_110_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_110_MPORT_238_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_110_MPORT_238_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_111_MPORT_111_en & tensorFile_111_MPORT_111_mask) begin
      tensorFile_111[tensorFile_111_MPORT_111_addr] <= tensorFile_111_MPORT_111_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_111_MPORT_239_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_111_MPORT_239_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_112_MPORT_112_en & tensorFile_112_MPORT_112_mask) begin
      tensorFile_112[tensorFile_112_MPORT_112_addr] <= tensorFile_112_MPORT_112_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_112_MPORT_240_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_112_MPORT_240_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_113_MPORT_113_en & tensorFile_113_MPORT_113_mask) begin
      tensorFile_113[tensorFile_113_MPORT_113_addr] <= tensorFile_113_MPORT_113_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_113_MPORT_241_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_113_MPORT_241_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_114_MPORT_114_en & tensorFile_114_MPORT_114_mask) begin
      tensorFile_114[tensorFile_114_MPORT_114_addr] <= tensorFile_114_MPORT_114_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_114_MPORT_242_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_114_MPORT_242_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_115_MPORT_115_en & tensorFile_115_MPORT_115_mask) begin
      tensorFile_115[tensorFile_115_MPORT_115_addr] <= tensorFile_115_MPORT_115_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_115_MPORT_243_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_115_MPORT_243_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_116_MPORT_116_en & tensorFile_116_MPORT_116_mask) begin
      tensorFile_116[tensorFile_116_MPORT_116_addr] <= tensorFile_116_MPORT_116_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_116_MPORT_244_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_116_MPORT_244_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_117_MPORT_117_en & tensorFile_117_MPORT_117_mask) begin
      tensorFile_117[tensorFile_117_MPORT_117_addr] <= tensorFile_117_MPORT_117_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_117_MPORT_245_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_117_MPORT_245_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_118_MPORT_118_en & tensorFile_118_MPORT_118_mask) begin
      tensorFile_118[tensorFile_118_MPORT_118_addr] <= tensorFile_118_MPORT_118_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_118_MPORT_246_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_118_MPORT_246_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_119_MPORT_119_en & tensorFile_119_MPORT_119_mask) begin
      tensorFile_119[tensorFile_119_MPORT_119_addr] <= tensorFile_119_MPORT_119_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_119_MPORT_247_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_119_MPORT_247_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_120_MPORT_120_en & tensorFile_120_MPORT_120_mask) begin
      tensorFile_120[tensorFile_120_MPORT_120_addr] <= tensorFile_120_MPORT_120_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_120_MPORT_248_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_120_MPORT_248_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_121_MPORT_121_en & tensorFile_121_MPORT_121_mask) begin
      tensorFile_121[tensorFile_121_MPORT_121_addr] <= tensorFile_121_MPORT_121_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_121_MPORT_249_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_121_MPORT_249_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_122_MPORT_122_en & tensorFile_122_MPORT_122_mask) begin
      tensorFile_122[tensorFile_122_MPORT_122_addr] <= tensorFile_122_MPORT_122_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_122_MPORT_250_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_122_MPORT_250_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_123_MPORT_123_en & tensorFile_123_MPORT_123_mask) begin
      tensorFile_123[tensorFile_123_MPORT_123_addr] <= tensorFile_123_MPORT_123_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_123_MPORT_251_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_123_MPORT_251_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_124_MPORT_124_en & tensorFile_124_MPORT_124_mask) begin
      tensorFile_124[tensorFile_124_MPORT_124_addr] <= tensorFile_124_MPORT_124_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_124_MPORT_252_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_124_MPORT_252_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_125_MPORT_125_en & tensorFile_125_MPORT_125_mask) begin
      tensorFile_125[tensorFile_125_MPORT_125_addr] <= tensorFile_125_MPORT_125_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_125_MPORT_253_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_125_MPORT_253_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_126_MPORT_126_en & tensorFile_126_MPORT_126_mask) begin
      tensorFile_126[tensorFile_126_MPORT_126_addr] <= tensorFile_126_MPORT_126_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_126_MPORT_254_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_126_MPORT_254_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if(tensorFile_127_MPORT_127_en & tensorFile_127_MPORT_127_mask) begin
      tensorFile_127[tensorFile_127_MPORT_127_addr] <= tensorFile_127_MPORT_127_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_127_MPORT_255_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_127_MPORT_255_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (reset) begin // @[TensorLoadNarrowVME.scala 54:22]
      state <= 1'h0; // @[TensorLoadNarrowVME.scala 54:22]
    end else begin
      state <= _GEN_1;
    end
    if (io_start) begin // @[TensorLoadNarrowVME.scala 88:18]
      blocksInFlight <= 17'h0; // @[TensorLoadNarrowVME.scala 89:20]
    end else if (state & _T & ~vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 90:66]
      blocksInFlight <= _blocksInFlight_T_1; // @[TensorLoadNarrowVME.scala 91:20]
    end else if (_T_1 & vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 92:65]
      blocksInFlight <= _blocksInFlight_T_5; // @[TensorLoadNarrowVME.scala 93:20]
    end else if (state & ~_T & vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 94:66]
      blocksInFlight <= _blocksInFlight_T_7; // @[TensorLoadNarrowVME.scala 96:20]
    end
    vmeDataBitsPipe_data <= io_vme_rd_data_bits_data; // @[TensorLoadNarrowVME.scala 67:32]
    vmeDataBitsPipe_tag <= io_vme_rd_data_bits_tag; // @[TensorLoadNarrowVME.scala 67:32]
    if (reset) begin // @[TensorLoadNarrowVME.scala 68:33]
      vmeDataValidPipe <= 1'h0; // @[TensorLoadNarrowVME.scala 68:33]
    end else begin
      vmeDataValidPipe <= io_vme_rd_data_valid; // @[TensorLoadNarrowVME.scala 68:33]
    end
    if (reset) begin // @[TensorLoadNarrowVME.scala 69:33]
      vmeDataReadyPipe <= 1'h0; // @[TensorLoadNarrowVME.scala 69:33]
    end else begin
      vmeDataReadyPipe <= io_vme_rd_data_ready; // @[TensorLoadNarrowVME.scala 69:33]
    end
    fillPadding_io_inst_REG <= io_inst; // @[TensorLoadNarrowVME.scala 121:33]
    if (reset) begin // @[TensorLoadNarrowVME.scala 122:34]
      fillPadding_io_start_REG <= 1'h0; // @[TensorLoadNarrowVME.scala 122:34]
    end else begin
      fillPadding_io_start_REG <= io_start; // @[TensorLoadNarrowVME.scala 122:34]
    end
    if (reset) begin // @[Reg.scala 27:20]
      rvalid <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      rvalid <= io_tensor_rd_0_idx_valid;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~io_start & ~_T_3 & ~_T_6 & _T_10 & ~(blocksInFlight > 17'h0 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorLoadNarrowVME.scala:95 assert(blocksInFlight > 0.U)\n"); // @[TensorLoadNarrowVME.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~io_start & ~_T_3 & ~_T_6 & _T_10 & ~(blocksInFlight > 17'h0 | reset)) begin
          $fatal; // @[TensorLoadNarrowVME.scala 95:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_0[initvar] = _RAND_0[63:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_1[initvar] = _RAND_3[63:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_2[initvar] = _RAND_6[63:0];
  _RAND_9 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_3[initvar] = _RAND_9[63:0];
  _RAND_12 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_4[initvar] = _RAND_12[63:0];
  _RAND_15 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_5[initvar] = _RAND_15[63:0];
  _RAND_18 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_6[initvar] = _RAND_18[63:0];
  _RAND_21 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_7[initvar] = _RAND_21[63:0];
  _RAND_24 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_8[initvar] = _RAND_24[63:0];
  _RAND_27 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_9[initvar] = _RAND_27[63:0];
  _RAND_30 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_10[initvar] = _RAND_30[63:0];
  _RAND_33 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_11[initvar] = _RAND_33[63:0];
  _RAND_36 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_12[initvar] = _RAND_36[63:0];
  _RAND_39 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_13[initvar] = _RAND_39[63:0];
  _RAND_42 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_14[initvar] = _RAND_42[63:0];
  _RAND_45 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_15[initvar] = _RAND_45[63:0];
  _RAND_48 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_16[initvar] = _RAND_48[63:0];
  _RAND_51 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_17[initvar] = _RAND_51[63:0];
  _RAND_54 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_18[initvar] = _RAND_54[63:0];
  _RAND_57 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_19[initvar] = _RAND_57[63:0];
  _RAND_60 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_20[initvar] = _RAND_60[63:0];
  _RAND_63 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_21[initvar] = _RAND_63[63:0];
  _RAND_66 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_22[initvar] = _RAND_66[63:0];
  _RAND_69 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_23[initvar] = _RAND_69[63:0];
  _RAND_72 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_24[initvar] = _RAND_72[63:0];
  _RAND_75 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_25[initvar] = _RAND_75[63:0];
  _RAND_78 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_26[initvar] = _RAND_78[63:0];
  _RAND_81 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_27[initvar] = _RAND_81[63:0];
  _RAND_84 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_28[initvar] = _RAND_84[63:0];
  _RAND_87 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_29[initvar] = _RAND_87[63:0];
  _RAND_90 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_30[initvar] = _RAND_90[63:0];
  _RAND_93 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_31[initvar] = _RAND_93[63:0];
  _RAND_96 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_32[initvar] = _RAND_96[63:0];
  _RAND_99 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_33[initvar] = _RAND_99[63:0];
  _RAND_102 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_34[initvar] = _RAND_102[63:0];
  _RAND_105 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_35[initvar] = _RAND_105[63:0];
  _RAND_108 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_36[initvar] = _RAND_108[63:0];
  _RAND_111 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_37[initvar] = _RAND_111[63:0];
  _RAND_114 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_38[initvar] = _RAND_114[63:0];
  _RAND_117 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_39[initvar] = _RAND_117[63:0];
  _RAND_120 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_40[initvar] = _RAND_120[63:0];
  _RAND_123 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_41[initvar] = _RAND_123[63:0];
  _RAND_126 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_42[initvar] = _RAND_126[63:0];
  _RAND_129 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_43[initvar] = _RAND_129[63:0];
  _RAND_132 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_44[initvar] = _RAND_132[63:0];
  _RAND_135 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_45[initvar] = _RAND_135[63:0];
  _RAND_138 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_46[initvar] = _RAND_138[63:0];
  _RAND_141 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_47[initvar] = _RAND_141[63:0];
  _RAND_144 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_48[initvar] = _RAND_144[63:0];
  _RAND_147 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_49[initvar] = _RAND_147[63:0];
  _RAND_150 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_50[initvar] = _RAND_150[63:0];
  _RAND_153 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_51[initvar] = _RAND_153[63:0];
  _RAND_156 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_52[initvar] = _RAND_156[63:0];
  _RAND_159 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_53[initvar] = _RAND_159[63:0];
  _RAND_162 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_54[initvar] = _RAND_162[63:0];
  _RAND_165 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_55[initvar] = _RAND_165[63:0];
  _RAND_168 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_56[initvar] = _RAND_168[63:0];
  _RAND_171 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_57[initvar] = _RAND_171[63:0];
  _RAND_174 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_58[initvar] = _RAND_174[63:0];
  _RAND_177 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_59[initvar] = _RAND_177[63:0];
  _RAND_180 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_60[initvar] = _RAND_180[63:0];
  _RAND_183 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_61[initvar] = _RAND_183[63:0];
  _RAND_186 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_62[initvar] = _RAND_186[63:0];
  _RAND_189 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_63[initvar] = _RAND_189[63:0];
  _RAND_192 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_64[initvar] = _RAND_192[63:0];
  _RAND_195 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_65[initvar] = _RAND_195[63:0];
  _RAND_198 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_66[initvar] = _RAND_198[63:0];
  _RAND_201 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_67[initvar] = _RAND_201[63:0];
  _RAND_204 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_68[initvar] = _RAND_204[63:0];
  _RAND_207 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_69[initvar] = _RAND_207[63:0];
  _RAND_210 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_70[initvar] = _RAND_210[63:0];
  _RAND_213 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_71[initvar] = _RAND_213[63:0];
  _RAND_216 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_72[initvar] = _RAND_216[63:0];
  _RAND_219 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_73[initvar] = _RAND_219[63:0];
  _RAND_222 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_74[initvar] = _RAND_222[63:0];
  _RAND_225 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_75[initvar] = _RAND_225[63:0];
  _RAND_228 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_76[initvar] = _RAND_228[63:0];
  _RAND_231 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_77[initvar] = _RAND_231[63:0];
  _RAND_234 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_78[initvar] = _RAND_234[63:0];
  _RAND_237 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_79[initvar] = _RAND_237[63:0];
  _RAND_240 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_80[initvar] = _RAND_240[63:0];
  _RAND_243 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_81[initvar] = _RAND_243[63:0];
  _RAND_246 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_82[initvar] = _RAND_246[63:0];
  _RAND_249 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_83[initvar] = _RAND_249[63:0];
  _RAND_252 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_84[initvar] = _RAND_252[63:0];
  _RAND_255 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_85[initvar] = _RAND_255[63:0];
  _RAND_258 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_86[initvar] = _RAND_258[63:0];
  _RAND_261 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_87[initvar] = _RAND_261[63:0];
  _RAND_264 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_88[initvar] = _RAND_264[63:0];
  _RAND_267 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_89[initvar] = _RAND_267[63:0];
  _RAND_270 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_90[initvar] = _RAND_270[63:0];
  _RAND_273 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_91[initvar] = _RAND_273[63:0];
  _RAND_276 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_92[initvar] = _RAND_276[63:0];
  _RAND_279 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_93[initvar] = _RAND_279[63:0];
  _RAND_282 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_94[initvar] = _RAND_282[63:0];
  _RAND_285 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_95[initvar] = _RAND_285[63:0];
  _RAND_288 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_96[initvar] = _RAND_288[63:0];
  _RAND_291 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_97[initvar] = _RAND_291[63:0];
  _RAND_294 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_98[initvar] = _RAND_294[63:0];
  _RAND_297 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_99[initvar] = _RAND_297[63:0];
  _RAND_300 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_100[initvar] = _RAND_300[63:0];
  _RAND_303 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_101[initvar] = _RAND_303[63:0];
  _RAND_306 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_102[initvar] = _RAND_306[63:0];
  _RAND_309 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_103[initvar] = _RAND_309[63:0];
  _RAND_312 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_104[initvar] = _RAND_312[63:0];
  _RAND_315 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_105[initvar] = _RAND_315[63:0];
  _RAND_318 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_106[initvar] = _RAND_318[63:0];
  _RAND_321 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_107[initvar] = _RAND_321[63:0];
  _RAND_324 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_108[initvar] = _RAND_324[63:0];
  _RAND_327 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_109[initvar] = _RAND_327[63:0];
  _RAND_330 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_110[initvar] = _RAND_330[63:0];
  _RAND_333 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_111[initvar] = _RAND_333[63:0];
  _RAND_336 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_112[initvar] = _RAND_336[63:0];
  _RAND_339 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_113[initvar] = _RAND_339[63:0];
  _RAND_342 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_114[initvar] = _RAND_342[63:0];
  _RAND_345 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_115[initvar] = _RAND_345[63:0];
  _RAND_348 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_116[initvar] = _RAND_348[63:0];
  _RAND_351 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_117[initvar] = _RAND_351[63:0];
  _RAND_354 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_118[initvar] = _RAND_354[63:0];
  _RAND_357 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_119[initvar] = _RAND_357[63:0];
  _RAND_360 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_120[initvar] = _RAND_360[63:0];
  _RAND_363 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_121[initvar] = _RAND_363[63:0];
  _RAND_366 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_122[initvar] = _RAND_366[63:0];
  _RAND_369 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_123[initvar] = _RAND_369[63:0];
  _RAND_372 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_124[initvar] = _RAND_372[63:0];
  _RAND_375 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_125[initvar] = _RAND_375[63:0];
  _RAND_378 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_126[initvar] = _RAND_378[63:0];
  _RAND_381 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    tensorFile_127[initvar] = _RAND_381[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tensorFile_0_MPORT_128_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tensorFile_0_MPORT_128_addr_pipe_0 = _RAND_2[9:0];
  _RAND_4 = {1{`RANDOM}};
  tensorFile_1_MPORT_129_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tensorFile_1_MPORT_129_addr_pipe_0 = _RAND_5[9:0];
  _RAND_7 = {1{`RANDOM}};
  tensorFile_2_MPORT_130_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tensorFile_2_MPORT_130_addr_pipe_0 = _RAND_8[9:0];
  _RAND_10 = {1{`RANDOM}};
  tensorFile_3_MPORT_131_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  tensorFile_3_MPORT_131_addr_pipe_0 = _RAND_11[9:0];
  _RAND_13 = {1{`RANDOM}};
  tensorFile_4_MPORT_132_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  tensorFile_4_MPORT_132_addr_pipe_0 = _RAND_14[9:0];
  _RAND_16 = {1{`RANDOM}};
  tensorFile_5_MPORT_133_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  tensorFile_5_MPORT_133_addr_pipe_0 = _RAND_17[9:0];
  _RAND_19 = {1{`RANDOM}};
  tensorFile_6_MPORT_134_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  tensorFile_6_MPORT_134_addr_pipe_0 = _RAND_20[9:0];
  _RAND_22 = {1{`RANDOM}};
  tensorFile_7_MPORT_135_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  tensorFile_7_MPORT_135_addr_pipe_0 = _RAND_23[9:0];
  _RAND_25 = {1{`RANDOM}};
  tensorFile_8_MPORT_136_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  tensorFile_8_MPORT_136_addr_pipe_0 = _RAND_26[9:0];
  _RAND_28 = {1{`RANDOM}};
  tensorFile_9_MPORT_137_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  tensorFile_9_MPORT_137_addr_pipe_0 = _RAND_29[9:0];
  _RAND_31 = {1{`RANDOM}};
  tensorFile_10_MPORT_138_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  tensorFile_10_MPORT_138_addr_pipe_0 = _RAND_32[9:0];
  _RAND_34 = {1{`RANDOM}};
  tensorFile_11_MPORT_139_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  tensorFile_11_MPORT_139_addr_pipe_0 = _RAND_35[9:0];
  _RAND_37 = {1{`RANDOM}};
  tensorFile_12_MPORT_140_en_pipe_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  tensorFile_12_MPORT_140_addr_pipe_0 = _RAND_38[9:0];
  _RAND_40 = {1{`RANDOM}};
  tensorFile_13_MPORT_141_en_pipe_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  tensorFile_13_MPORT_141_addr_pipe_0 = _RAND_41[9:0];
  _RAND_43 = {1{`RANDOM}};
  tensorFile_14_MPORT_142_en_pipe_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  tensorFile_14_MPORT_142_addr_pipe_0 = _RAND_44[9:0];
  _RAND_46 = {1{`RANDOM}};
  tensorFile_15_MPORT_143_en_pipe_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  tensorFile_15_MPORT_143_addr_pipe_0 = _RAND_47[9:0];
  _RAND_49 = {1{`RANDOM}};
  tensorFile_16_MPORT_144_en_pipe_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  tensorFile_16_MPORT_144_addr_pipe_0 = _RAND_50[9:0];
  _RAND_52 = {1{`RANDOM}};
  tensorFile_17_MPORT_145_en_pipe_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  tensorFile_17_MPORT_145_addr_pipe_0 = _RAND_53[9:0];
  _RAND_55 = {1{`RANDOM}};
  tensorFile_18_MPORT_146_en_pipe_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  tensorFile_18_MPORT_146_addr_pipe_0 = _RAND_56[9:0];
  _RAND_58 = {1{`RANDOM}};
  tensorFile_19_MPORT_147_en_pipe_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  tensorFile_19_MPORT_147_addr_pipe_0 = _RAND_59[9:0];
  _RAND_61 = {1{`RANDOM}};
  tensorFile_20_MPORT_148_en_pipe_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  tensorFile_20_MPORT_148_addr_pipe_0 = _RAND_62[9:0];
  _RAND_64 = {1{`RANDOM}};
  tensorFile_21_MPORT_149_en_pipe_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tensorFile_21_MPORT_149_addr_pipe_0 = _RAND_65[9:0];
  _RAND_67 = {1{`RANDOM}};
  tensorFile_22_MPORT_150_en_pipe_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  tensorFile_22_MPORT_150_addr_pipe_0 = _RAND_68[9:0];
  _RAND_70 = {1{`RANDOM}};
  tensorFile_23_MPORT_151_en_pipe_0 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  tensorFile_23_MPORT_151_addr_pipe_0 = _RAND_71[9:0];
  _RAND_73 = {1{`RANDOM}};
  tensorFile_24_MPORT_152_en_pipe_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  tensorFile_24_MPORT_152_addr_pipe_0 = _RAND_74[9:0];
  _RAND_76 = {1{`RANDOM}};
  tensorFile_25_MPORT_153_en_pipe_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  tensorFile_25_MPORT_153_addr_pipe_0 = _RAND_77[9:0];
  _RAND_79 = {1{`RANDOM}};
  tensorFile_26_MPORT_154_en_pipe_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  tensorFile_26_MPORT_154_addr_pipe_0 = _RAND_80[9:0];
  _RAND_82 = {1{`RANDOM}};
  tensorFile_27_MPORT_155_en_pipe_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  tensorFile_27_MPORT_155_addr_pipe_0 = _RAND_83[9:0];
  _RAND_85 = {1{`RANDOM}};
  tensorFile_28_MPORT_156_en_pipe_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  tensorFile_28_MPORT_156_addr_pipe_0 = _RAND_86[9:0];
  _RAND_88 = {1{`RANDOM}};
  tensorFile_29_MPORT_157_en_pipe_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  tensorFile_29_MPORT_157_addr_pipe_0 = _RAND_89[9:0];
  _RAND_91 = {1{`RANDOM}};
  tensorFile_30_MPORT_158_en_pipe_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  tensorFile_30_MPORT_158_addr_pipe_0 = _RAND_92[9:0];
  _RAND_94 = {1{`RANDOM}};
  tensorFile_31_MPORT_159_en_pipe_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  tensorFile_31_MPORT_159_addr_pipe_0 = _RAND_95[9:0];
  _RAND_97 = {1{`RANDOM}};
  tensorFile_32_MPORT_160_en_pipe_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  tensorFile_32_MPORT_160_addr_pipe_0 = _RAND_98[9:0];
  _RAND_100 = {1{`RANDOM}};
  tensorFile_33_MPORT_161_en_pipe_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  tensorFile_33_MPORT_161_addr_pipe_0 = _RAND_101[9:0];
  _RAND_103 = {1{`RANDOM}};
  tensorFile_34_MPORT_162_en_pipe_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  tensorFile_34_MPORT_162_addr_pipe_0 = _RAND_104[9:0];
  _RAND_106 = {1{`RANDOM}};
  tensorFile_35_MPORT_163_en_pipe_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  tensorFile_35_MPORT_163_addr_pipe_0 = _RAND_107[9:0];
  _RAND_109 = {1{`RANDOM}};
  tensorFile_36_MPORT_164_en_pipe_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  tensorFile_36_MPORT_164_addr_pipe_0 = _RAND_110[9:0];
  _RAND_112 = {1{`RANDOM}};
  tensorFile_37_MPORT_165_en_pipe_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  tensorFile_37_MPORT_165_addr_pipe_0 = _RAND_113[9:0];
  _RAND_115 = {1{`RANDOM}};
  tensorFile_38_MPORT_166_en_pipe_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  tensorFile_38_MPORT_166_addr_pipe_0 = _RAND_116[9:0];
  _RAND_118 = {1{`RANDOM}};
  tensorFile_39_MPORT_167_en_pipe_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  tensorFile_39_MPORT_167_addr_pipe_0 = _RAND_119[9:0];
  _RAND_121 = {1{`RANDOM}};
  tensorFile_40_MPORT_168_en_pipe_0 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  tensorFile_40_MPORT_168_addr_pipe_0 = _RAND_122[9:0];
  _RAND_124 = {1{`RANDOM}};
  tensorFile_41_MPORT_169_en_pipe_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  tensorFile_41_MPORT_169_addr_pipe_0 = _RAND_125[9:0];
  _RAND_127 = {1{`RANDOM}};
  tensorFile_42_MPORT_170_en_pipe_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  tensorFile_42_MPORT_170_addr_pipe_0 = _RAND_128[9:0];
  _RAND_130 = {1{`RANDOM}};
  tensorFile_43_MPORT_171_en_pipe_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  tensorFile_43_MPORT_171_addr_pipe_0 = _RAND_131[9:0];
  _RAND_133 = {1{`RANDOM}};
  tensorFile_44_MPORT_172_en_pipe_0 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  tensorFile_44_MPORT_172_addr_pipe_0 = _RAND_134[9:0];
  _RAND_136 = {1{`RANDOM}};
  tensorFile_45_MPORT_173_en_pipe_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  tensorFile_45_MPORT_173_addr_pipe_0 = _RAND_137[9:0];
  _RAND_139 = {1{`RANDOM}};
  tensorFile_46_MPORT_174_en_pipe_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  tensorFile_46_MPORT_174_addr_pipe_0 = _RAND_140[9:0];
  _RAND_142 = {1{`RANDOM}};
  tensorFile_47_MPORT_175_en_pipe_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  tensorFile_47_MPORT_175_addr_pipe_0 = _RAND_143[9:0];
  _RAND_145 = {1{`RANDOM}};
  tensorFile_48_MPORT_176_en_pipe_0 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  tensorFile_48_MPORT_176_addr_pipe_0 = _RAND_146[9:0];
  _RAND_148 = {1{`RANDOM}};
  tensorFile_49_MPORT_177_en_pipe_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  tensorFile_49_MPORT_177_addr_pipe_0 = _RAND_149[9:0];
  _RAND_151 = {1{`RANDOM}};
  tensorFile_50_MPORT_178_en_pipe_0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  tensorFile_50_MPORT_178_addr_pipe_0 = _RAND_152[9:0];
  _RAND_154 = {1{`RANDOM}};
  tensorFile_51_MPORT_179_en_pipe_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  tensorFile_51_MPORT_179_addr_pipe_0 = _RAND_155[9:0];
  _RAND_157 = {1{`RANDOM}};
  tensorFile_52_MPORT_180_en_pipe_0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  tensorFile_52_MPORT_180_addr_pipe_0 = _RAND_158[9:0];
  _RAND_160 = {1{`RANDOM}};
  tensorFile_53_MPORT_181_en_pipe_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  tensorFile_53_MPORT_181_addr_pipe_0 = _RAND_161[9:0];
  _RAND_163 = {1{`RANDOM}};
  tensorFile_54_MPORT_182_en_pipe_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  tensorFile_54_MPORT_182_addr_pipe_0 = _RAND_164[9:0];
  _RAND_166 = {1{`RANDOM}};
  tensorFile_55_MPORT_183_en_pipe_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  tensorFile_55_MPORT_183_addr_pipe_0 = _RAND_167[9:0];
  _RAND_169 = {1{`RANDOM}};
  tensorFile_56_MPORT_184_en_pipe_0 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  tensorFile_56_MPORT_184_addr_pipe_0 = _RAND_170[9:0];
  _RAND_172 = {1{`RANDOM}};
  tensorFile_57_MPORT_185_en_pipe_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  tensorFile_57_MPORT_185_addr_pipe_0 = _RAND_173[9:0];
  _RAND_175 = {1{`RANDOM}};
  tensorFile_58_MPORT_186_en_pipe_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  tensorFile_58_MPORT_186_addr_pipe_0 = _RAND_176[9:0];
  _RAND_178 = {1{`RANDOM}};
  tensorFile_59_MPORT_187_en_pipe_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  tensorFile_59_MPORT_187_addr_pipe_0 = _RAND_179[9:0];
  _RAND_181 = {1{`RANDOM}};
  tensorFile_60_MPORT_188_en_pipe_0 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  tensorFile_60_MPORT_188_addr_pipe_0 = _RAND_182[9:0];
  _RAND_184 = {1{`RANDOM}};
  tensorFile_61_MPORT_189_en_pipe_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  tensorFile_61_MPORT_189_addr_pipe_0 = _RAND_185[9:0];
  _RAND_187 = {1{`RANDOM}};
  tensorFile_62_MPORT_190_en_pipe_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  tensorFile_62_MPORT_190_addr_pipe_0 = _RAND_188[9:0];
  _RAND_190 = {1{`RANDOM}};
  tensorFile_63_MPORT_191_en_pipe_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  tensorFile_63_MPORT_191_addr_pipe_0 = _RAND_191[9:0];
  _RAND_193 = {1{`RANDOM}};
  tensorFile_64_MPORT_192_en_pipe_0 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  tensorFile_64_MPORT_192_addr_pipe_0 = _RAND_194[9:0];
  _RAND_196 = {1{`RANDOM}};
  tensorFile_65_MPORT_193_en_pipe_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  tensorFile_65_MPORT_193_addr_pipe_0 = _RAND_197[9:0];
  _RAND_199 = {1{`RANDOM}};
  tensorFile_66_MPORT_194_en_pipe_0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  tensorFile_66_MPORT_194_addr_pipe_0 = _RAND_200[9:0];
  _RAND_202 = {1{`RANDOM}};
  tensorFile_67_MPORT_195_en_pipe_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  tensorFile_67_MPORT_195_addr_pipe_0 = _RAND_203[9:0];
  _RAND_205 = {1{`RANDOM}};
  tensorFile_68_MPORT_196_en_pipe_0 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  tensorFile_68_MPORT_196_addr_pipe_0 = _RAND_206[9:0];
  _RAND_208 = {1{`RANDOM}};
  tensorFile_69_MPORT_197_en_pipe_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  tensorFile_69_MPORT_197_addr_pipe_0 = _RAND_209[9:0];
  _RAND_211 = {1{`RANDOM}};
  tensorFile_70_MPORT_198_en_pipe_0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  tensorFile_70_MPORT_198_addr_pipe_0 = _RAND_212[9:0];
  _RAND_214 = {1{`RANDOM}};
  tensorFile_71_MPORT_199_en_pipe_0 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  tensorFile_71_MPORT_199_addr_pipe_0 = _RAND_215[9:0];
  _RAND_217 = {1{`RANDOM}};
  tensorFile_72_MPORT_200_en_pipe_0 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  tensorFile_72_MPORT_200_addr_pipe_0 = _RAND_218[9:0];
  _RAND_220 = {1{`RANDOM}};
  tensorFile_73_MPORT_201_en_pipe_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  tensorFile_73_MPORT_201_addr_pipe_0 = _RAND_221[9:0];
  _RAND_223 = {1{`RANDOM}};
  tensorFile_74_MPORT_202_en_pipe_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  tensorFile_74_MPORT_202_addr_pipe_0 = _RAND_224[9:0];
  _RAND_226 = {1{`RANDOM}};
  tensorFile_75_MPORT_203_en_pipe_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  tensorFile_75_MPORT_203_addr_pipe_0 = _RAND_227[9:0];
  _RAND_229 = {1{`RANDOM}};
  tensorFile_76_MPORT_204_en_pipe_0 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  tensorFile_76_MPORT_204_addr_pipe_0 = _RAND_230[9:0];
  _RAND_232 = {1{`RANDOM}};
  tensorFile_77_MPORT_205_en_pipe_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  tensorFile_77_MPORT_205_addr_pipe_0 = _RAND_233[9:0];
  _RAND_235 = {1{`RANDOM}};
  tensorFile_78_MPORT_206_en_pipe_0 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  tensorFile_78_MPORT_206_addr_pipe_0 = _RAND_236[9:0];
  _RAND_238 = {1{`RANDOM}};
  tensorFile_79_MPORT_207_en_pipe_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  tensorFile_79_MPORT_207_addr_pipe_0 = _RAND_239[9:0];
  _RAND_241 = {1{`RANDOM}};
  tensorFile_80_MPORT_208_en_pipe_0 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  tensorFile_80_MPORT_208_addr_pipe_0 = _RAND_242[9:0];
  _RAND_244 = {1{`RANDOM}};
  tensorFile_81_MPORT_209_en_pipe_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  tensorFile_81_MPORT_209_addr_pipe_0 = _RAND_245[9:0];
  _RAND_247 = {1{`RANDOM}};
  tensorFile_82_MPORT_210_en_pipe_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  tensorFile_82_MPORT_210_addr_pipe_0 = _RAND_248[9:0];
  _RAND_250 = {1{`RANDOM}};
  tensorFile_83_MPORT_211_en_pipe_0 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  tensorFile_83_MPORT_211_addr_pipe_0 = _RAND_251[9:0];
  _RAND_253 = {1{`RANDOM}};
  tensorFile_84_MPORT_212_en_pipe_0 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  tensorFile_84_MPORT_212_addr_pipe_0 = _RAND_254[9:0];
  _RAND_256 = {1{`RANDOM}};
  tensorFile_85_MPORT_213_en_pipe_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  tensorFile_85_MPORT_213_addr_pipe_0 = _RAND_257[9:0];
  _RAND_259 = {1{`RANDOM}};
  tensorFile_86_MPORT_214_en_pipe_0 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  tensorFile_86_MPORT_214_addr_pipe_0 = _RAND_260[9:0];
  _RAND_262 = {1{`RANDOM}};
  tensorFile_87_MPORT_215_en_pipe_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  tensorFile_87_MPORT_215_addr_pipe_0 = _RAND_263[9:0];
  _RAND_265 = {1{`RANDOM}};
  tensorFile_88_MPORT_216_en_pipe_0 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  tensorFile_88_MPORT_216_addr_pipe_0 = _RAND_266[9:0];
  _RAND_268 = {1{`RANDOM}};
  tensorFile_89_MPORT_217_en_pipe_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  tensorFile_89_MPORT_217_addr_pipe_0 = _RAND_269[9:0];
  _RAND_271 = {1{`RANDOM}};
  tensorFile_90_MPORT_218_en_pipe_0 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  tensorFile_90_MPORT_218_addr_pipe_0 = _RAND_272[9:0];
  _RAND_274 = {1{`RANDOM}};
  tensorFile_91_MPORT_219_en_pipe_0 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  tensorFile_91_MPORT_219_addr_pipe_0 = _RAND_275[9:0];
  _RAND_277 = {1{`RANDOM}};
  tensorFile_92_MPORT_220_en_pipe_0 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  tensorFile_92_MPORT_220_addr_pipe_0 = _RAND_278[9:0];
  _RAND_280 = {1{`RANDOM}};
  tensorFile_93_MPORT_221_en_pipe_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  tensorFile_93_MPORT_221_addr_pipe_0 = _RAND_281[9:0];
  _RAND_283 = {1{`RANDOM}};
  tensorFile_94_MPORT_222_en_pipe_0 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  tensorFile_94_MPORT_222_addr_pipe_0 = _RAND_284[9:0];
  _RAND_286 = {1{`RANDOM}};
  tensorFile_95_MPORT_223_en_pipe_0 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  tensorFile_95_MPORT_223_addr_pipe_0 = _RAND_287[9:0];
  _RAND_289 = {1{`RANDOM}};
  tensorFile_96_MPORT_224_en_pipe_0 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  tensorFile_96_MPORT_224_addr_pipe_0 = _RAND_290[9:0];
  _RAND_292 = {1{`RANDOM}};
  tensorFile_97_MPORT_225_en_pipe_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  tensorFile_97_MPORT_225_addr_pipe_0 = _RAND_293[9:0];
  _RAND_295 = {1{`RANDOM}};
  tensorFile_98_MPORT_226_en_pipe_0 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  tensorFile_98_MPORT_226_addr_pipe_0 = _RAND_296[9:0];
  _RAND_298 = {1{`RANDOM}};
  tensorFile_99_MPORT_227_en_pipe_0 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  tensorFile_99_MPORT_227_addr_pipe_0 = _RAND_299[9:0];
  _RAND_301 = {1{`RANDOM}};
  tensorFile_100_MPORT_228_en_pipe_0 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  tensorFile_100_MPORT_228_addr_pipe_0 = _RAND_302[9:0];
  _RAND_304 = {1{`RANDOM}};
  tensorFile_101_MPORT_229_en_pipe_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  tensorFile_101_MPORT_229_addr_pipe_0 = _RAND_305[9:0];
  _RAND_307 = {1{`RANDOM}};
  tensorFile_102_MPORT_230_en_pipe_0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  tensorFile_102_MPORT_230_addr_pipe_0 = _RAND_308[9:0];
  _RAND_310 = {1{`RANDOM}};
  tensorFile_103_MPORT_231_en_pipe_0 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  tensorFile_103_MPORT_231_addr_pipe_0 = _RAND_311[9:0];
  _RAND_313 = {1{`RANDOM}};
  tensorFile_104_MPORT_232_en_pipe_0 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  tensorFile_104_MPORT_232_addr_pipe_0 = _RAND_314[9:0];
  _RAND_316 = {1{`RANDOM}};
  tensorFile_105_MPORT_233_en_pipe_0 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  tensorFile_105_MPORT_233_addr_pipe_0 = _RAND_317[9:0];
  _RAND_319 = {1{`RANDOM}};
  tensorFile_106_MPORT_234_en_pipe_0 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  tensorFile_106_MPORT_234_addr_pipe_0 = _RAND_320[9:0];
  _RAND_322 = {1{`RANDOM}};
  tensorFile_107_MPORT_235_en_pipe_0 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  tensorFile_107_MPORT_235_addr_pipe_0 = _RAND_323[9:0];
  _RAND_325 = {1{`RANDOM}};
  tensorFile_108_MPORT_236_en_pipe_0 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  tensorFile_108_MPORT_236_addr_pipe_0 = _RAND_326[9:0];
  _RAND_328 = {1{`RANDOM}};
  tensorFile_109_MPORT_237_en_pipe_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  tensorFile_109_MPORT_237_addr_pipe_0 = _RAND_329[9:0];
  _RAND_331 = {1{`RANDOM}};
  tensorFile_110_MPORT_238_en_pipe_0 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  tensorFile_110_MPORT_238_addr_pipe_0 = _RAND_332[9:0];
  _RAND_334 = {1{`RANDOM}};
  tensorFile_111_MPORT_239_en_pipe_0 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  tensorFile_111_MPORT_239_addr_pipe_0 = _RAND_335[9:0];
  _RAND_337 = {1{`RANDOM}};
  tensorFile_112_MPORT_240_en_pipe_0 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  tensorFile_112_MPORT_240_addr_pipe_0 = _RAND_338[9:0];
  _RAND_340 = {1{`RANDOM}};
  tensorFile_113_MPORT_241_en_pipe_0 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  tensorFile_113_MPORT_241_addr_pipe_0 = _RAND_341[9:0];
  _RAND_343 = {1{`RANDOM}};
  tensorFile_114_MPORT_242_en_pipe_0 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  tensorFile_114_MPORT_242_addr_pipe_0 = _RAND_344[9:0];
  _RAND_346 = {1{`RANDOM}};
  tensorFile_115_MPORT_243_en_pipe_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  tensorFile_115_MPORT_243_addr_pipe_0 = _RAND_347[9:0];
  _RAND_349 = {1{`RANDOM}};
  tensorFile_116_MPORT_244_en_pipe_0 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  tensorFile_116_MPORT_244_addr_pipe_0 = _RAND_350[9:0];
  _RAND_352 = {1{`RANDOM}};
  tensorFile_117_MPORT_245_en_pipe_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  tensorFile_117_MPORT_245_addr_pipe_0 = _RAND_353[9:0];
  _RAND_355 = {1{`RANDOM}};
  tensorFile_118_MPORT_246_en_pipe_0 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  tensorFile_118_MPORT_246_addr_pipe_0 = _RAND_356[9:0];
  _RAND_358 = {1{`RANDOM}};
  tensorFile_119_MPORT_247_en_pipe_0 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  tensorFile_119_MPORT_247_addr_pipe_0 = _RAND_359[9:0];
  _RAND_361 = {1{`RANDOM}};
  tensorFile_120_MPORT_248_en_pipe_0 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  tensorFile_120_MPORT_248_addr_pipe_0 = _RAND_362[9:0];
  _RAND_364 = {1{`RANDOM}};
  tensorFile_121_MPORT_249_en_pipe_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  tensorFile_121_MPORT_249_addr_pipe_0 = _RAND_365[9:0];
  _RAND_367 = {1{`RANDOM}};
  tensorFile_122_MPORT_250_en_pipe_0 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  tensorFile_122_MPORT_250_addr_pipe_0 = _RAND_368[9:0];
  _RAND_370 = {1{`RANDOM}};
  tensorFile_123_MPORT_251_en_pipe_0 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  tensorFile_123_MPORT_251_addr_pipe_0 = _RAND_371[9:0];
  _RAND_373 = {1{`RANDOM}};
  tensorFile_124_MPORT_252_en_pipe_0 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  tensorFile_124_MPORT_252_addr_pipe_0 = _RAND_374[9:0];
  _RAND_376 = {1{`RANDOM}};
  tensorFile_125_MPORT_253_en_pipe_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  tensorFile_125_MPORT_253_addr_pipe_0 = _RAND_377[9:0];
  _RAND_379 = {1{`RANDOM}};
  tensorFile_126_MPORT_254_en_pipe_0 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  tensorFile_126_MPORT_254_addr_pipe_0 = _RAND_380[9:0];
  _RAND_382 = {1{`RANDOM}};
  tensorFile_127_MPORT_255_en_pipe_0 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  tensorFile_127_MPORT_255_addr_pipe_0 = _RAND_383[9:0];
  _RAND_384 = {1{`RANDOM}};
  state = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  blocksInFlight = _RAND_385[16:0];
  _RAND_386 = {2{`RANDOM}};
  vmeDataBitsPipe_data = _RAND_386[63:0];
  _RAND_387 = {1{`RANDOM}};
  vmeDataBitsPipe_tag = _RAND_387[20:0];
  _RAND_388 = {1{`RANDOM}};
  vmeDataValidPipe = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  vmeDataReadyPipe = _RAND_389[0:0];
  _RAND_390 = {4{`RANDOM}};
  fillPadding_io_inst_REG = _RAND_390[127:0];
  _RAND_391 = {1{`RANDOM}};
  fillPadding_io_start_REG = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  rvalid = _RAND_392[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule