module Pipe(
  input   clock,
  input   reset,
  input   io_enq_valid,
  input   io_enq_bits,
  output  io_deq_valid,
  output  io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  io_deq_v; // @[Valid.scala 117:22]
  reg  io_deq_b; // @[Reg.scala 15:16]
  reg  io_deq_outPipe_valid; // @[Valid.scala 117:22]
  reg  io_deq_outPipe_bits; // @[Reg.scala 15:16]
  reg  io_deq_outPipe_valid_1; // @[Valid.scala 117:22]
  reg  io_deq_outPipe_bits_1; // @[Reg.scala 15:16]
  assign io_deq_valid = io_deq_outPipe_valid_1; // @[Valid.scala 112:21 Valid.scala 113:17]
  assign io_deq_bits = io_deq_outPipe_bits_1; // @[Valid.scala 112:21 Valid.scala 114:16]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 117:22]
      io_deq_v <= 1'h0; // @[Valid.scala 117:22]
    end else begin
      io_deq_v <= io_enq_valid; // @[Valid.scala 117:22]
    end
    if (io_enq_valid) begin // @[Reg.scala 16:19]
      io_deq_b <= io_enq_bits; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Valid.scala 117:22]
      io_deq_outPipe_valid <= 1'h0; // @[Valid.scala 117:22]
    end else begin
      io_deq_outPipe_valid <= io_deq_v; // @[Valid.scala 117:22]
    end
    if (io_deq_v) begin // @[Reg.scala 16:19]
      io_deq_outPipe_bits <= io_deq_b; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Valid.scala 117:22]
      io_deq_outPipe_valid_1 <= 1'h0; // @[Valid.scala 117:22]
    end else begin
      io_deq_outPipe_valid_1 <= io_deq_outPipe_valid; // @[Valid.scala 117:22]
    end
    if (io_deq_outPipe_valid) begin // @[Reg.scala 16:19]
      io_deq_outPipe_bits_1 <= io_deq_outPipe_bits; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_deq_v = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_deq_b = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_deq_outPipe_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  io_deq_outPipe_bits = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_deq_outPipe_valid_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_deq_outPipe_bits_1 = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule